LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE IEEE.std_logic_misc.all;
USE work.typeDeclarations.all;

ENTITY audioROM IS
PORT(
	clk: in std_logic;
	audio_request: in std_logic;
	keys: in std_logic_vector (15 downto 0);
	octave: in std_logic_vector (1 downto 0);
	z: out unsigned (15 downto 0)
);
END ENTITY audioROM;

ARCHITECTURE rom OF audioROM IS

COMPONENT SampleAdder16 IS
PORT(
		keys: in std_logic_vector(15 downto 0);

		a: in unsigned(15 downto 0);
		b: in unsigned(15 downto 0);
		c: in unsigned(15 downto 0);
		d: in unsigned(15 downto 0);
		e: in unsigned(15 downto 0);
		f: in unsigned(15 downto 0);
		g: in unsigned(15 downto 0);
		h: in unsigned(15 downto 0);
		i: in unsigned(15 downto 0);
		j: in unsigned(15 downto 0);
		k: in unsigned(15 downto 0);
		l: in unsigned(15 downto 0);
		m: in unsigned(15 downto 0);
		n: in unsigned(15 downto 0);
		o: in unsigned(15 downto 0);
		p: in unsigned(15 downto 0);
		
		z: out unsigned(15 downto 0)
);
END COMPONENT SampleAdder16;

COMPONENT SampleContainer IS
PORT(
		clk: in std_logic;
		stream: in std_logic;
		rom1, rom2, rom3: in hex;
		loop1, loop2, loop3: in natural;
		octave: in std_logic_vector (1 downto 0);
		audio_request: in std_logic;
		z: out unsigned (15 downto 0)
);
END COMPONENT SampleContainer;

SIGNAL k0, k1, k2, k3, k4, k5, k6, k7, k8, k9, k10, k11, k12, k13, k14, k15: unsigned (15 downto 0) := X"0000";

CONSTANT num_samples: nat_num := (
	--indexing set by octave(1) - tone(2)
	000 => 103,
	001 => 109,
	002 => 116,
	003 => 123,
	004 => 130,
	005 => 138,
	006 => 147,
	007 => 155,
	008 => 165,
	009 => 174,
	010 => 185,
	011 => 196,
	012 => 207,
	013 => 220,
	014 => 233,
	015 => 247,
	100 => 51,
	101 => 54,
	102 => 58,
	103 => 61,
	104 => 65,
	105 => 69,
	106 => 73,
	107 => 77,
	108 => 82,
	109 => 87,
	110 => 92,
	111 => 97,
	112 => 103,
	113 => 109,
	114 => 116,
	115 => 123,
	200 => 51,
	201 => 54,
	202 => 58,
	203 => 61,
	204 => 25,
	205 => 27,
	206 => 28,
	207 => 30,
	208 => 32,
	209 => 34,
	210 => 36,
	211 => 38,
	212 => 41,
	213 => 43,
	214 => 46,
	215 => 48,
	others => 0
);

CONSTANT C3: hex := (
	000 => X"0000",
	001 => X"033E",
	002 => X"067B",
	003 => X"09B8",
	004 => X"0CF2",
	005 => X"102B",
	006 => X"1361",
	007 => X"1694",
	008 => X"19C3",
	009 => X"1CEE",
	010 => X"2015",
	011 => X"2336",
	012 => X"2651",
	013 => X"2966",
	014 => X"2C74",
	015 => X"2F7A",
	016 => X"3279",
	017 => X"3570",
	018 => X"385E",
	019 => X"3B43",
	020 => X"3E1D",
	021 => X"40EE",
	022 => X"43B4",
	023 => X"466F",
	024 => X"491E",
	025 => X"4BC2",
	026 => X"4E58",
	027 => X"50E2",
	028 => X"535F",
	029 => X"55CE",
	030 => X"582F",
	031 => X"5A81",
	032 => X"5CC5",
	033 => X"5EF9",
	034 => X"611E",
	035 => X"6332",
	036 => X"6537",
	037 => X"672B",
	038 => X"690D",
	039 => X"6ADF",
	040 => X"6C9F",
	041 => X"6E4D",
	042 => X"6FE9",
	043 => X"7173",
	044 => X"72EA",
	045 => X"744E",
	046 => X"759F",
	047 => X"76DD",
	048 => X"7807",
	049 => X"791D",
	050 => X"7A20",
	051 => X"7B0E",
	052 => X"7BE8",
	053 => X"7CAE",
	054 => X"7D60",
	055 => X"7DFD",
	056 => X"7E85",
	057 => X"7EF8",
	058 => X"7F56",
	059 => X"7FA0",
	060 => X"7FD4",
	061 => X"7FF4",
	062 => X"7FFF",
	063 => X"7FF4",
	064 => X"7FD4",
	065 => X"7FA0",
	066 => X"7F56",
	067 => X"7EF8",
	068 => X"7E85",
	069 => X"7DFD",
	070 => X"7D60",
	071 => X"7CAE",
	072 => X"7BE8",
	073 => X"7B0E",
	074 => X"7A20",
	075 => X"791D",
	076 => X"7807",
	077 => X"76DD",
	078 => X"759F",
	079 => X"744E",
	080 => X"72EA",
	081 => X"7173",
	082 => X"6FE9",
	083 => X"6E4D",
	084 => X"6C9F",
	085 => X"6ADF",
	086 => X"690D",
	087 => X"672B",
	088 => X"6537",
	089 => X"6332",
	090 => X"611E",
	091 => X"5EF9",
	092 => X"5CC5",
	093 => X"5A81",
	094 => X"582F",
	095 => X"55CE",
	096 => X"535F",
	097 => X"50E2",
	098 => X"4E58",
	099 => X"4BC2",
	100 => X"491E",
	101 => X"466F",
	102 => X"43B4",
	103 => X"40EE",
	104 => X"3E1D",
	105 => X"3B43",
	106 => X"385E",
	107 => X"3570",
	108 => X"3279",
	109 => X"2F7A",
	110 => X"2C74",
	111 => X"2966",
	112 => X"2651",
	113 => X"2336",
	114 => X"2015",
	115 => X"1CEE",
	116 => X"19C3",
	117 => X"1694",
	118 => X"1361",
	119 => X"102B",
	120 => X"0CF2",
	121 => X"09B8",
	122 => X"067B",
	123 => X"033E",
	124 => X"0000",
	125 => X"FCC0",
	126 => X"F983",
	127 => X"F646",
	128 => X"F30C",
	129 => X"EFD3",
	130 => X"EC9D",
	131 => X"E96A",
	132 => X"E63B",
	133 => X"E310",
	134 => X"DFE9",
	135 => X"DCC8",
	136 => X"D9AD",
	137 => X"D698",
	138 => X"D38A",
	139 => X"D084",
	140 => X"CD85",
	141 => X"CA8E",
	142 => X"C7A0",
	143 => X"C4BB",
	144 => X"C1E1",
	145 => X"BF10",
	146 => X"BC4A",
	147 => X"B98F",
	148 => X"B6E0",
	149 => X"B43C",
	150 => X"B1A6",
	151 => X"AF1C",
	152 => X"AC9F",
	153 => X"AA30",
	154 => X"A7CF",
	155 => X"A57D",
	156 => X"A339",
	157 => X"A105",
	158 => X"9EE0",
	159 => X"9CCC",
	160 => X"9AC7",
	161 => X"98D3",
	162 => X"96F1",
	163 => X"951F",
	164 => X"935F",
	165 => X"91B1",
	166 => X"9015",
	167 => X"8E8B",
	168 => X"8D14",
	169 => X"8BB0",
	170 => X"8A5F",
	171 => X"8921",
	172 => X"87F7",
	173 => X"86E1",
	174 => X"85DE",
	175 => X"84F0",
	176 => X"8416",
	177 => X"8350",
	178 => X"829E",
	179 => X"8201",
	180 => X"8179",
	181 => X"8106",
	182 => X"80A8",
	183 => X"805E",
	184 => X"802A",
	185 => X"800A",
	186 => X"8000",
	187 => X"800A",
	188 => X"802A",
	189 => X"805E",
	190 => X"80A8",
	191 => X"8106",
	192 => X"8179",
	193 => X"8201",
	194 => X"829E",
	195 => X"8350",
	196 => X"8416",
	197 => X"84F0",
	198 => X"85DE",
	199 => X"86E1",
	200 => X"87F7",
	201 => X"8921",
	202 => X"8A5F",
	203 => X"8BB0",
	204 => X"8D14",
	205 => X"8E8B",
	206 => X"9015",
	207 => X"91B1",
	208 => X"935F",
	209 => X"951F",
	210 => X"96F1",
	211 => X"98D3",
	212 => X"9AC7",
	213 => X"9CCC",
	214 => X"9EE0",
	215 => X"A105",
	216 => X"A339",
	217 => X"A57D",
	218 => X"A7CF",
	219 => X"AA30",
	220 => X"AC9F",
	221 => X"AF1C",
	222 => X"B1A6",
	223 => X"B43C",
	224 => X"B6E0",
	225 => X"B98F",
	226 => X"BC4A",
	227 => X"BF10",
	228 => X"C1E1",
	229 => X"C4BB",
	230 => X"C7A0",
	231 => X"CA8E",
	232 => X"CD85",
	233 => X"D084",
	234 => X"D38A",
	235 => X"D698",
	236 => X"D9AD",
	237 => X"DCC8",
	238 => X"DFE9",
	239 => X"E310",
	240 => X"E63B",
	241 => X"E96A",
	242 => X"EC9D",
	243 => X"EFD3",
	244 => X"F30C",
	245 => X"F646",
	246 => X"F983",
	247 => X"FCC0",
	others => X"0000"
);

CONSTANT CS3: hex := (
	000 => X"0000",
	001 => X"036F",
	002 => X"06DE",
	003 => X"0A4C",
	004 => X"0DB8",
	005 => X"1121",
	006 => X"1488",
	007 => X"17EA",
	008 => X"1B48",
	009 => X"1EA1",
	010 => X"21F4",
	011 => X"2542",
	012 => X"2888",
	013 => X"2BC6",
	014 => X"2EFD",
	015 => X"322B",
	016 => X"3550",
	017 => X"386B",
	018 => X"3B7B",
	019 => X"3E81",
	020 => X"417A",
	021 => X"4468",
	022 => X"474A",
	023 => X"4A1E",
	024 => X"4CE4",
	025 => X"4F9C",
	026 => X"5246",
	027 => X"54E0",
	028 => X"576B",
	029 => X"59E5",
	030 => X"5C4F",
	031 => X"5EA8",
	032 => X"60EF",
	033 => X"6325",
	034 => X"6548",
	035 => X"6759",
	036 => X"6956",
	037 => X"6B40",
	038 => X"6D16",
	039 => X"6ED9",
	040 => X"7086",
	041 => X"721F",
	042 => X"73A3",
	043 => X"7511",
	044 => X"766A",
	045 => X"77AD",
	046 => X"78DA",
	047 => X"79F1",
	048 => X"7AF1",
	049 => X"7BDA",
	050 => X"7CAD",
	051 => X"7D68",
	052 => X"7E0D",
	053 => X"7E9A",
	054 => X"7F10",
	055 => X"7F6E",
	056 => X"7FB5",
	057 => X"7FE4",
	058 => X"7FFC",
	059 => X"7FFC",
	060 => X"7FE4",
	061 => X"7FB5",
	062 => X"7F6E",
	063 => X"7F10",
	064 => X"7E9A",
	065 => X"7E0D",
	066 => X"7D68",
	067 => X"7CAD",
	068 => X"7BDA",
	069 => X"7AF1",
	070 => X"79F1",
	071 => X"78DA",
	072 => X"77AD",
	073 => X"766A",
	074 => X"7511",
	075 => X"73A3",
	076 => X"721F",
	077 => X"7086",
	078 => X"6ED9",
	079 => X"6D16",
	080 => X"6B40",
	081 => X"6956",
	082 => X"6759",
	083 => X"6548",
	084 => X"6325",
	085 => X"60EF",
	086 => X"5EA8",
	087 => X"5C4F",
	088 => X"59E5",
	089 => X"576B",
	090 => X"54E0",
	091 => X"5246",
	092 => X"4F9C",
	093 => X"4CE4",
	094 => X"4A1E",
	095 => X"474A",
	096 => X"4468",
	097 => X"417A",
	098 => X"3E81",
	099 => X"3B7B",
	100 => X"386B",
	101 => X"3550",
	102 => X"322B",
	103 => X"2EFD",
	104 => X"2BC6",
	105 => X"2888",
	106 => X"2542",
	107 => X"21F4",
	108 => X"1EA1",
	109 => X"1B48",
	110 => X"17EA",
	111 => X"1488",
	112 => X"1121",
	113 => X"0DB8",
	114 => X"0A4C",
	115 => X"06DE",
	116 => X"036F",
	117 => X"FFFE",
	118 => X"FC8F",
	119 => X"F920",
	120 => X"F5B2",
	121 => X"F246",
	122 => X"EEDD",
	123 => X"EB76",
	124 => X"E814",
	125 => X"E4B6",
	126 => X"E15D",
	127 => X"DE0A",
	128 => X"DABC",
	129 => X"D776",
	130 => X"D438",
	131 => X"D101",
	132 => X"CDD3",
	133 => X"CAAE",
	134 => X"C793",
	135 => X"C483",
	136 => X"C17D",
	137 => X"BE84",
	138 => X"BB96",
	139 => X"B8B4",
	140 => X"B5E0",
	141 => X"B31A",
	142 => X"B062",
	143 => X"ADB8",
	144 => X"AB1E",
	145 => X"A893",
	146 => X"A619",
	147 => X"A3AF",
	148 => X"A156",
	149 => X"9F0F",
	150 => X"9CD9",
	151 => X"9AB6",
	152 => X"98A5",
	153 => X"96A8",
	154 => X"94BE",
	155 => X"92E8",
	156 => X"9125",
	157 => X"8F78",
	158 => X"8DDF",
	159 => X"8C5B",
	160 => X"8AED",
	161 => X"8994",
	162 => X"8851",
	163 => X"8724",
	164 => X"860D",
	165 => X"850D",
	166 => X"8424",
	167 => X"8351",
	168 => X"8296",
	169 => X"81F1",
	170 => X"8164",
	171 => X"80EE",
	172 => X"8090",
	173 => X"8049",
	174 => X"801A",
	175 => X"8002",
	176 => X"8002",
	177 => X"801A",
	178 => X"8049",
	179 => X"8090",
	180 => X"80EE",
	181 => X"8164",
	182 => X"81F1",
	183 => X"8296",
	184 => X"8351",
	185 => X"8424",
	186 => X"850D",
	187 => X"860D",
	188 => X"8724",
	189 => X"8851",
	190 => X"8994",
	191 => X"8AED",
	192 => X"8C5B",
	193 => X"8DDF",
	194 => X"8F78",
	195 => X"9125",
	196 => X"92E8",
	197 => X"94BE",
	198 => X"96A8",
	199 => X"98A5",
	200 => X"9AB6",
	201 => X"9CD9",
	202 => X"9F0F",
	203 => X"A156",
	204 => X"A3AF",
	205 => X"A619",
	206 => X"A893",
	207 => X"AB1E",
	208 => X"ADB8",
	209 => X"B062",
	210 => X"B31A",
	211 => X"B5E0",
	212 => X"B8B4",
	213 => X"BB96",
	214 => X"BE84",
	215 => X"C17D",
	216 => X"C483",
	217 => X"C793",
	218 => X"CAAE",
	219 => X"CDD3",
	220 => X"D101",
	221 => X"D438",
	222 => X"D776",
	223 => X"DABC",
	224 => X"DE0A",
	225 => X"E15D",
	226 => X"E4B6",
	227 => X"E814",
	228 => X"EB76",
	229 => X"EEDD",
	230 => X"F246",
	231 => X"F5B2",
	232 => X"F920",
	233 => X"FC8F",
	234 => X"0000",
	235 => X"036F",
	236 => X"06DE",
	237 => X"0A4C",
	238 => X"0DB8",
	239 => X"1121",
	240 => X"1488",
	241 => X"17EA",
	242 => X"1B48",
	243 => X"1EA1",
	244 => X"21F4",
	245 => X"2542",
	246 => X"2888",
	247 => X"2BC6",
	others => X"0000"
);

CONSTANT D3: hex := (
	000 => X"0000",
	001 => X"03A3",
	002 => X"0746",
	003 => X"0AE7",
	004 => X"0E86",
	005 => X"1222",
	006 => X"15BA",
	007 => X"194E",
	008 => X"1CDC",
	009 => X"2065",
	010 => X"23E6",
	011 => X"2761",
	012 => X"2AD3",
	013 => X"2E3C",
	014 => X"319C",
	015 => X"34F2",
	016 => X"383C",
	017 => X"3B7B",
	018 => X"3EAE",
	019 => X"41D3",
	020 => X"44EB",
	021 => X"47F5",
	022 => X"4AF0",
	023 => X"4DDB",
	024 => X"50B7",
	025 => X"5381",
	026 => X"563A",
	027 => X"58E2",
	028 => X"5B77",
	029 => X"5DF9",
	030 => X"6068",
	031 => X"62C2",
	032 => X"6509",
	033 => X"673A",
	034 => X"6956",
	035 => X"6B5C",
	036 => X"6D4C",
	037 => X"6F26",
	038 => X"70E8",
	039 => X"7293",
	040 => X"7427",
	041 => X"75A2",
	042 => X"7705",
	043 => X"784F",
	044 => X"7981",
	045 => X"7A99",
	046 => X"7B98",
	047 => X"7C7D",
	048 => X"7D49",
	049 => X"7DFB",
	050 => X"7E92",
	051 => X"7F10",
	052 => X"7F73",
	053 => X"7FBB",
	054 => X"7FEA",
	055 => X"7FFE",
	056 => X"7FF7",
	057 => X"7FD6",
	058 => X"7F9A",
	059 => X"7F44",
	060 => X"7ED4",
	061 => X"7E4A",
	062 => X"7DA5",
	063 => X"7CE6",
	064 => X"7C0E",
	065 => X"7B1C",
	066 => X"7A10",
	067 => X"78EB",
	068 => X"77AD",
	069 => X"7656",
	070 => X"74E7",
	071 => X"7360",
	072 => X"71C1",
	073 => X"700A",
	074 => X"6E3C",
	075 => X"6C57",
	076 => X"6A5C",
	077 => X"684B",
	078 => X"6624",
	079 => X"63E8",
	080 => X"6198",
	081 => X"5F33",
	082 => X"5CBA",
	083 => X"5A2F",
	084 => X"5790",
	085 => X"54E0",
	086 => X"521E",
	087 => X"4F4B",
	088 => X"4C68",
	089 => X"4974",
	090 => X"4672",
	091 => X"4361",
	092 => X"4042",
	093 => X"3D16",
	094 => X"39DD",
	095 => X"3698",
	096 => X"3348",
	097 => X"2FED",
	098 => X"2C89",
	099 => X"291B",
	100 => X"25A5",
	101 => X"2226",
	102 => X"1EA1",
	103 => X"1B16",
	104 => X"1784",
	105 => X"13EE",
	106 => X"1054",
	107 => X"0CB7",
	108 => X"0917",
	109 => X"0574",
	110 => X"01D1",
	111 => X"FE2D",
	112 => X"FA8A",
	113 => X"F6E7",
	114 => X"F347",
	115 => X"EFAA",
	116 => X"EC10",
	117 => X"E87A",
	118 => X"E4E8",
	119 => X"E15D",
	120 => X"DDD8",
	121 => X"DA59",
	122 => X"D6E3",
	123 => X"D375",
	124 => X"D011",
	125 => X"CCB6",
	126 => X"C966",
	127 => X"C621",
	128 => X"C2E8",
	129 => X"BFBC",
	130 => X"BC9D",
	131 => X"B98C",
	132 => X"B68A",
	133 => X"B396",
	134 => X"B0B3",
	135 => X"ADE0",
	136 => X"AB1E",
	137 => X"A86E",
	138 => X"A5CF",
	139 => X"A344",
	140 => X"A0CB",
	141 => X"9E66",
	142 => X"9C16",
	143 => X"99DA",
	144 => X"97B3",
	145 => X"95A2",
	146 => X"93A7",
	147 => X"91C2",
	148 => X"8FF4",
	149 => X"8E3D",
	150 => X"8C9E",
	151 => X"8B17",
	152 => X"89A8",
	153 => X"8851",
	154 => X"8713",
	155 => X"85EE",
	156 => X"84E2",
	157 => X"83F0",
	158 => X"8318",
	159 => X"8259",
	160 => X"81B4",
	161 => X"812A",
	162 => X"80BA",
	163 => X"8064",
	164 => X"8028",
	165 => X"8007",
	166 => X"8000",
	167 => X"8014",
	168 => X"8043",
	169 => X"808B",
	170 => X"80EE",
	171 => X"816C",
	172 => X"8203",
	173 => X"82B5",
	174 => X"8381",
	175 => X"8466",
	176 => X"8565",
	177 => X"867D",
	178 => X"87AF",
	179 => X"88F9",
	180 => X"8A5C",
	181 => X"8BD7",
	182 => X"8D6B",
	183 => X"8F16",
	184 => X"90D8",
	185 => X"92B2",
	186 => X"94A2",
	187 => X"96A8",
	188 => X"98C4",
	189 => X"9AF5",
	190 => X"9D3C",
	191 => X"9F96",
	192 => X"A205",
	193 => X"A487",
	194 => X"A71C",
	195 => X"A9C4",
	196 => X"AC7D",
	197 => X"AF47",
	198 => X"B223",
	199 => X"B50E",
	200 => X"B809",
	201 => X"BB13",
	202 => X"BE2B",
	203 => X"C150",
	204 => X"C483",
	205 => X"C7C2",
	206 => X"CB0C",
	207 => X"CE62",
	208 => X"D1C2",
	209 => X"D52B",
	210 => X"D89D",
	211 => X"DC18",
	212 => X"DF99",
	213 => X"E322",
	214 => X"E6B0",
	215 => X"EA44",
	216 => X"EDDC",
	217 => X"F178",
	218 => X"F517",
	219 => X"F8B8",
	220 => X"FC5B",
	221 => X"0000",
	222 => X"03A3",
	223 => X"0746",
	224 => X"0AE7",
	225 => X"0E86",
	226 => X"1222",
	227 => X"15BA",
	228 => X"194E",
	229 => X"1CDC",
	230 => X"2065",
	231 => X"23E6",
	232 => X"2761",
	233 => X"2AD3",
	234 => X"2E3C",
	235 => X"319C",
	236 => X"34F2",
	237 => X"383C",
	238 => X"3B7B",
	239 => X"3EAE",
	240 => X"41D3",
	241 => X"44EB",
	242 => X"47F5",
	243 => X"4AF0",
	244 => X"4DDB",
	245 => X"50B7",
	246 => X"5381",
	247 => X"563A",
	others => X"0000"
);

CONSTANT DS3: hex := (
	000 => X"0000",
	001 => X"03DD",
	002 => X"07BA",
	003 => X"0B95",
	004 => X"0F6D",
	005 => X"1342",
	006 => X"1712",
	007 => X"1ADD",
	008 => X"1EA1",
	009 => X"225E",
	010 => X"2614",
	011 => X"29C0",
	012 => X"2D63",
	013 => X"30FB",
	014 => X"3487",
	015 => X"3808",
	016 => X"3B7B",
	017 => X"3EE0",
	018 => X"4237",
	019 => X"457E",
	020 => X"48B5",
	021 => X"4BDB",
	022 => X"4EF0",
	023 => X"51F1",
	024 => X"54E0",
	025 => X"57BB",
	026 => X"5A81",
	027 => X"5D32",
	028 => X"5FCE",
	029 => X"6253",
	030 => X"64C1",
	031 => X"6718",
	032 => X"6956",
	033 => X"6B7C",
	034 => X"6D89",
	035 => X"6F7C",
	036 => X"7155",
	037 => X"7314",
	038 => X"74B8",
	039 => X"7640",
	040 => X"77AD",
	041 => X"78FE",
	042 => X"7A33",
	043 => X"7B4B",
	044 => X"7C46",
	045 => X"7D25",
	046 => X"7DE6",
	047 => X"7E89",
	048 => X"7F10",
	049 => X"7F78",
	050 => X"7FC3",
	051 => X"7FF0",
	052 => X"7FFF",
	053 => X"7FF0",
	054 => X"7FC3",
	055 => X"7F78",
	056 => X"7F10",
	057 => X"7E89",
	058 => X"7DE6",
	059 => X"7D25",
	060 => X"7C46",
	061 => X"7B4B",
	062 => X"7A33",
	063 => X"78FE",
	064 => X"77AD",
	065 => X"7640",
	066 => X"74B8",
	067 => X"7314",
	068 => X"7155",
	069 => X"6F7C",
	070 => X"6D89",
	071 => X"6B7C",
	072 => X"6956",
	073 => X"6718",
	074 => X"64C1",
	075 => X"6253",
	076 => X"5FCE",
	077 => X"5D32",
	078 => X"5A81",
	079 => X"57BB",
	080 => X"54E0",
	081 => X"51F1",
	082 => X"4EF0",
	083 => X"4BDB",
	084 => X"48B5",
	085 => X"457E",
	086 => X"4237",
	087 => X"3EE0",
	088 => X"3B7B",
	089 => X"3808",
	090 => X"3487",
	091 => X"30FB",
	092 => X"2D63",
	093 => X"29C0",
	094 => X"2614",
	095 => X"225E",
	096 => X"1EA1",
	097 => X"1ADD",
	098 => X"1712",
	099 => X"1342",
	100 => X"0F6D",
	101 => X"0B95",
	102 => X"07BA",
	103 => X"03DD",
	104 => X"0000",
	105 => X"FC21",
	106 => X"F844",
	107 => X"F469",
	108 => X"F091",
	109 => X"ECBC",
	110 => X"E8EC",
	111 => X"E521",
	112 => X"E15D",
	113 => X"DDA0",
	114 => X"D9EA",
	115 => X"D63E",
	116 => X"D29B",
	117 => X"CF03",
	118 => X"CB77",
	119 => X"C7F6",
	120 => X"C483",
	121 => X"C11E",
	122 => X"BDC7",
	123 => X"BA80",
	124 => X"B749",
	125 => X"B423",
	126 => X"B10E",
	127 => X"AE0D",
	128 => X"AB1E",
	129 => X"A843",
	130 => X"A57D",
	131 => X"A2CC",
	132 => X"A030",
	133 => X"9DAB",
	134 => X"9B3D",
	135 => X"98E6",
	136 => X"96A8",
	137 => X"9482",
	138 => X"9275",
	139 => X"9082",
	140 => X"8EA9",
	141 => X"8CEA",
	142 => X"8B46",
	143 => X"89BE",
	144 => X"8851",
	145 => X"8700",
	146 => X"85CB",
	147 => X"84B3",
	148 => X"83B8",
	149 => X"82D9",
	150 => X"8218",
	151 => X"8175",
	152 => X"80EE",
	153 => X"8086",
	154 => X"803B",
	155 => X"800E",
	156 => X"8000",
	157 => X"800E",
	158 => X"803B",
	159 => X"8086",
	160 => X"80EE",
	161 => X"8175",
	162 => X"8218",
	163 => X"82D9",
	164 => X"83B8",
	165 => X"84B3",
	166 => X"85CB",
	167 => X"8700",
	168 => X"8851",
	169 => X"89BE",
	170 => X"8B46",
	171 => X"8CEA",
	172 => X"8EA9",
	173 => X"9082",
	174 => X"9275",
	175 => X"9482",
	176 => X"96A8",
	177 => X"98E6",
	178 => X"9B3D",
	179 => X"9DAB",
	180 => X"A030",
	181 => X"A2CC",
	182 => X"A57D",
	183 => X"A843",
	184 => X"AB1E",
	185 => X"AE0D",
	186 => X"B10E",
	187 => X"B423",
	188 => X"B749",
	189 => X"BA80",
	190 => X"BDC7",
	191 => X"C11E",
	192 => X"C483",
	193 => X"C7F6",
	194 => X"CB77",
	195 => X"CF03",
	196 => X"D29B",
	197 => X"D63E",
	198 => X"D9EA",
	199 => X"DDA0",
	200 => X"E15D",
	201 => X"E521",
	202 => X"E8EC",
	203 => X"ECBC",
	204 => X"F091",
	205 => X"F469",
	206 => X"F844",
	207 => X"FC21",
	208 => X"FFFE",
	209 => X"03DD",
	210 => X"07BA",
	211 => X"0B95",
	212 => X"0F6D",
	213 => X"1342",
	214 => X"1712",
	215 => X"1ADD",
	216 => X"1EA1",
	217 => X"225E",
	218 => X"2614",
	219 => X"29C0",
	220 => X"2D63",
	221 => X"30FB",
	222 => X"3487",
	223 => X"3808",
	224 => X"3B7B",
	225 => X"3EE0",
	226 => X"4237",
	227 => X"457E",
	228 => X"48B5",
	229 => X"4BDB",
	230 => X"4EF0",
	231 => X"51F1",
	232 => X"54E0",
	233 => X"57BB",
	234 => X"5A81",
	235 => X"5D32",
	236 => X"5FCE",
	237 => X"6253",
	238 => X"64C1",
	239 => X"6718",
	240 => X"6956",
	241 => X"6B7C",
	242 => X"6D89",
	243 => X"6F7C",
	244 => X"7155",
	245 => X"7314",
	246 => X"74B8",
	247 => X"7640",
	others => X"0000"
);

CONSTANT E3: hex := (
	000 => X"0000",
	001 => X"0414",
	002 => X"0828",
	003 => X"0C3A",
	004 => X"1048",
	005 => X"1453",
	006 => X"1858",
	007 => X"1C56",
	008 => X"204E",
	009 => X"243D",
	010 => X"2822",
	011 => X"2BFD",
	012 => X"2FCD",
	013 => X"3390",
	014 => X"3745",
	015 => X"3AED",
	016 => X"3E84",
	017 => X"420C",
	018 => X"4583",
	019 => X"48E7",
	020 => X"4C38",
	021 => X"4F76",
	022 => X"529F",
	023 => X"55B2",
	024 => X"58AF",
	025 => X"5B95",
	026 => X"5E63",
	027 => X"6118",
	028 => X"63B4",
	029 => X"6637",
	030 => X"689E",
	031 => X"6AEB",
	032 => X"6D1B",
	033 => X"6F2F",
	034 => X"7126",
	035 => X"7300",
	036 => X"74BC",
	037 => X"7659",
	038 => X"77D8",
	039 => X"7937",
	040 => X"7A77",
	041 => X"7B97",
	042 => X"7C96",
	043 => X"7D76",
	044 => X"7E34",
	045 => X"7ED2",
	046 => X"7F4F",
	047 => X"7FAA",
	048 => X"7FE4",
	049 => X"7FFD",
	050 => X"7FF5",
	051 => X"7FCB",
	052 => X"7F81",
	053 => X"7F14",
	054 => X"7E87",
	055 => X"7DD9",
	056 => X"7D0A",
	057 => X"7C1B",
	058 => X"7B0B",
	059 => X"79DB",
	060 => X"788B",
	061 => X"771C",
	062 => X"758E",
	063 => X"73E2",
	064 => X"7217",
	065 => X"702E",
	066 => X"6E29",
	067 => X"6C06",
	068 => X"69C8",
	069 => X"676E",
	070 => X"64F9",
	071 => X"626A",
	072 => X"5FC1",
	073 => X"5CFF",
	074 => X"5A25",
	075 => X"5733",
	076 => X"542B",
	077 => X"510D",
	078 => X"4DDA",
	079 => X"4A92",
	080 => X"4737",
	081 => X"43CA",
	082 => X"404A",
	083 => X"3CBA",
	084 => X"391B",
	085 => X"356C",
	086 => X"31B0",
	087 => X"2DE6",
	088 => X"2A11",
	089 => X"2631",
	090 => X"2246",
	091 => X"1E53",
	092 => X"1A58",
	093 => X"1656",
	094 => X"124E",
	095 => X"0E42",
	096 => X"0A31",
	097 => X"061F",
	098 => X"020A",
	099 => X"FDF4",
	100 => X"F9DF",
	101 => X"F5CD",
	102 => X"F1BC",
	103 => X"EDB0",
	104 => X"E9A8",
	105 => X"E5A6",
	106 => X"E1AB",
	107 => X"DDB8",
	108 => X"D9CD",
	109 => X"D5ED",
	110 => X"D218",
	111 => X"CE4E",
	112 => X"CA92",
	113 => X"C6E3",
	114 => X"C344",
	115 => X"BFB4",
	116 => X"BC34",
	117 => X"B8C7",
	118 => X"B56C",
	119 => X"B224",
	120 => X"AEF1",
	121 => X"ABD3",
	122 => X"A8CB",
	123 => X"A5D9",
	124 => X"A2FF",
	125 => X"A03D",
	126 => X"9D94",
	127 => X"9B05",
	128 => X"9890",
	129 => X"9636",
	130 => X"93F8",
	131 => X"91D5",
	132 => X"8FD0",
	133 => X"8DE7",
	134 => X"8C1C",
	135 => X"8A70",
	136 => X"88E2",
	137 => X"8773",
	138 => X"8623",
	139 => X"84F3",
	140 => X"83E3",
	141 => X"82F4",
	142 => X"8225",
	143 => X"8177",
	144 => X"80EA",
	145 => X"807D",
	146 => X"8033",
	147 => X"8009",
	148 => X"8001",
	149 => X"801A",
	150 => X"8054",
	151 => X"80AF",
	152 => X"812C",
	153 => X"81CA",
	154 => X"8288",
	155 => X"8368",
	156 => X"8467",
	157 => X"8587",
	158 => X"86C7",
	159 => X"8826",
	160 => X"89A5",
	161 => X"8B42",
	162 => X"8CFE",
	163 => X"8ED8",
	164 => X"90CF",
	165 => X"92E3",
	166 => X"9513",
	167 => X"9760",
	168 => X"99C7",
	169 => X"9C4A",
	170 => X"9EE6",
	171 => X"A19B",
	172 => X"A469",
	173 => X"A74F",
	174 => X"AA4C",
	175 => X"AD5F",
	176 => X"B088",
	177 => X"B3C6",
	178 => X"B717",
	179 => X"BA7B",
	180 => X"BDF2",
	181 => X"C17A",
	182 => X"C511",
	183 => X"C8B9",
	184 => X"CC6E",
	185 => X"D031",
	186 => X"D401",
	187 => X"D7DC",
	188 => X"DBC1",
	189 => X"DFB0",
	190 => X"E3A8",
	191 => X"E7A6",
	192 => X"EBAB",
	193 => X"EFB6",
	194 => X"F3C4",
	195 => X"F7D6",
	196 => X"FBEA",
	197 => X"0000",
	198 => X"0414",
	199 => X"0828",
	200 => X"0C3A",
	201 => X"1048",
	202 => X"1453",
	203 => X"1858",
	204 => X"1C56",
	205 => X"204E",
	206 => X"243D",
	207 => X"2822",
	208 => X"2BFD",
	209 => X"2FCD",
	210 => X"3390",
	211 => X"3745",
	212 => X"3AED",
	213 => X"3E84",
	214 => X"420C",
	215 => X"4583",
	216 => X"48E7",
	217 => X"4C38",
	218 => X"4F76",
	219 => X"529F",
	220 => X"55B2",
	221 => X"58AF",
	222 => X"5B95",
	223 => X"5E63",
	224 => X"6118",
	225 => X"63B4",
	226 => X"6637",
	227 => X"689E",
	228 => X"6AEB",
	229 => X"6D1B",
	230 => X"6F2F",
	231 => X"7126",
	232 => X"7300",
	233 => X"74BC",
	234 => X"7659",
	235 => X"77D8",
	236 => X"7937",
	237 => X"7A77",
	238 => X"7B97",
	239 => X"7C96",
	240 => X"7D76",
	241 => X"7E34",
	242 => X"7ED2",
	243 => X"7F4F",
	244 => X"7FAA",
	245 => X"7FE4",
	246 => X"7FFD",
	247 => X"7FF5",
	others => X"0000"
);

CONSTANT F3: hex := (
	000 => X"0000",
	001 => X"0452",
	002 => X"08A4",
	003 => X"0CF2",
	004 => X"113E",
	005 => X"1584",
	006 => X"19C3",
	007 => X"1DFC",
	008 => X"222B",
	009 => X"2651",
	010 => X"2A6B",
	011 => X"2E79",
	012 => X"3279",
	013 => X"366B",
	014 => X"3A4D",
	015 => X"3E1D",
	016 => X"41DC",
	017 => X"4587",
	018 => X"491E",
	019 => X"4CA0",
	020 => X"500B",
	021 => X"535F",
	022 => X"569B",
	023 => X"59BD",
	024 => X"5CC5",
	025 => X"5FB2",
	026 => X"6283",
	027 => X"6537",
	028 => X"67CD",
	029 => X"6A46",
	030 => X"6C9F",
	031 => X"6ED9",
	032 => X"70F2",
	033 => X"72EA",
	034 => X"74C0",
	035 => X"7675",
	036 => X"7807",
	037 => X"7976",
	038 => X"7AC1",
	039 => X"7BE8",
	040 => X"7CEC",
	041 => X"7DCB",
	042 => X"7E85",
	043 => X"7F1A",
	044 => X"7F8A",
	045 => X"7FD4",
	046 => X"7FFA",
	047 => X"7FFA",
	048 => X"7FD4",
	049 => X"7F8A",
	050 => X"7F1A",
	051 => X"7E85",
	052 => X"7DCB",
	053 => X"7CEC",
	054 => X"7BE8",
	055 => X"7AC1",
	056 => X"7976",
	057 => X"7807",
	058 => X"7675",
	059 => X"74C0",
	060 => X"72EA",
	061 => X"70F2",
	062 => X"6ED9",
	063 => X"6C9F",
	064 => X"6A46",
	065 => X"67CD",
	066 => X"6537",
	067 => X"6283",
	068 => X"5FB2",
	069 => X"5CC5",
	070 => X"59BD",
	071 => X"569B",
	072 => X"535F",
	073 => X"500B",
	074 => X"4CA0",
	075 => X"491E",
	076 => X"4587",
	077 => X"41DC",
	078 => X"3E1D",
	079 => X"3A4D",
	080 => X"366B",
	081 => X"3279",
	082 => X"2E79",
	083 => X"2A6B",
	084 => X"2651",
	085 => X"222B",
	086 => X"1DFC",
	087 => X"19C3",
	088 => X"1584",
	089 => X"113E",
	090 => X"0CF2",
	091 => X"08A4",
	092 => X"0452",
	093 => X"FFFE",
	094 => X"FBAC",
	095 => X"F75A",
	096 => X"F30C",
	097 => X"EEC0",
	098 => X"EA7A",
	099 => X"E63B",
	100 => X"E202",
	101 => X"DDD3",
	102 => X"D9AD",
	103 => X"D593",
	104 => X"D185",
	105 => X"CD85",
	106 => X"C993",
	107 => X"C5B1",
	108 => X"C1E1",
	109 => X"BE22",
	110 => X"BA77",
	111 => X"B6E0",
	112 => X"B35E",
	113 => X"AFF3",
	114 => X"AC9F",
	115 => X"A963",
	116 => X"A641",
	117 => X"A339",
	118 => X"A04C",
	119 => X"9D7B",
	120 => X"9AC7",
	121 => X"9831",
	122 => X"95B8",
	123 => X"935F",
	124 => X"9125",
	125 => X"8F0C",
	126 => X"8D14",
	127 => X"8B3E",
	128 => X"8989",
	129 => X"87F7",
	130 => X"8688",
	131 => X"853D",
	132 => X"8416",
	133 => X"8312",
	134 => X"8233",
	135 => X"8179",
	136 => X"80E4",
	137 => X"8074",
	138 => X"802A",
	139 => X"8004",
	140 => X"8004",
	141 => X"802A",
	142 => X"8074",
	143 => X"80E4",
	144 => X"8179",
	145 => X"8233",
	146 => X"8312",
	147 => X"8416",
	148 => X"853D",
	149 => X"8688",
	150 => X"87F7",
	151 => X"8989",
	152 => X"8B3E",
	153 => X"8D14",
	154 => X"8F0C",
	155 => X"9125",
	156 => X"935F",
	157 => X"95B8",
	158 => X"9831",
	159 => X"9AC7",
	160 => X"9D7B",
	161 => X"A04C",
	162 => X"A339",
	163 => X"A641",
	164 => X"A963",
	165 => X"AC9F",
	166 => X"AFF3",
	167 => X"B35E",
	168 => X"B6E0",
	169 => X"BA77",
	170 => X"BE22",
	171 => X"C1E1",
	172 => X"C5B1",
	173 => X"C993",
	174 => X"CD85",
	175 => X"D185",
	176 => X"D593",
	177 => X"D9AD",
	178 => X"DDD3",
	179 => X"E202",
	180 => X"E63B",
	181 => X"EA7A",
	182 => X"EEC0",
	183 => X"F30C",
	184 => X"F75A",
	185 => X"FBAC",
	186 => X"0000",
	187 => X"0452",
	188 => X"08A4",
	189 => X"0CF2",
	190 => X"113E",
	191 => X"1584",
	192 => X"19C3",
	193 => X"1DFC",
	194 => X"222B",
	195 => X"2651",
	196 => X"2A6B",
	197 => X"2E79",
	198 => X"3279",
	199 => X"366B",
	200 => X"3A4D",
	201 => X"3E1D",
	202 => X"41DC",
	203 => X"4587",
	204 => X"491E",
	205 => X"4CA0",
	206 => X"500B",
	207 => X"535F",
	208 => X"569B",
	209 => X"59BD",
	210 => X"5CC5",
	211 => X"5FB2",
	212 => X"6283",
	213 => X"6537",
	214 => X"67CD",
	215 => X"6A46",
	216 => X"6C9F",
	217 => X"6ED9",
	218 => X"70F2",
	219 => X"72EA",
	220 => X"74C0",
	221 => X"7675",
	222 => X"7807",
	223 => X"7976",
	224 => X"7AC1",
	225 => X"7BE8",
	226 => X"7CEC",
	227 => X"7DCB",
	228 => X"7E85",
	229 => X"7F1A",
	230 => X"7F8A",
	231 => X"7FD4",
	232 => X"7FFA",
	233 => X"7FFA",
	234 => X"7FD4",
	235 => X"7F8A",
	236 => X"7F1A",
	237 => X"7E85",
	238 => X"7DCB",
	239 => X"7CEC",
	240 => X"7BE8",
	241 => X"7AC1",
	242 => X"7976",
	243 => X"7807",
	244 => X"7675",
	245 => X"74C0",
	246 => X"72EA",
	247 => X"70F2",
	others => X"0000"
);

CONSTANT FS3: hex := (
	000 => X"0000",
	001 => X"0498",
	002 => X"092E",
	003 => X"0DC2",
	004 => X"1251",
	005 => X"16DA",
	006 => X"1B5C",
	007 => X"1FD4",
	008 => X"2442",
	009 => X"28A4",
	010 => X"2CF9",
	011 => X"313F",
	012 => X"3574",
	013 => X"3998",
	014 => X"3DA9",
	015 => X"41A6",
	016 => X"458D",
	017 => X"495C",
	018 => X"4D14",
	019 => X"50B3",
	020 => X"5436",
	021 => X"579E",
	022 => X"5AE9",
	023 => X"5E16",
	024 => X"6124",
	025 => X"6412",
	026 => X"66DF",
	027 => X"698A",
	028 => X"6C12",
	029 => X"6E76",
	030 => X"70B6",
	031 => X"72D1",
	032 => X"74C6",
	033 => X"7694",
	034 => X"783B",
	035 => X"79BB",
	036 => X"7B12",
	037 => X"7C41",
	038 => X"7D47",
	039 => X"7E23",
	040 => X"7ED6",
	041 => X"7F5F",
	042 => X"7FBE",
	043 => X"7FF3",
	044 => X"7FFD",
	045 => X"7FDE",
	046 => X"7F94",
	047 => X"7F20",
	048 => X"7E82",
	049 => X"7DBA",
	050 => X"7CC9",
	051 => X"7BAF",
	052 => X"7A6C",
	053 => X"7900",
	054 => X"776D",
	055 => X"75B2",
	056 => X"73D0",
	057 => X"71C8",
	058 => X"6F9B",
	059 => X"6D48",
	060 => X"6AD2",
	061 => X"6838",
	062 => X"657C",
	063 => X"629F",
	064 => X"5FA1",
	065 => X"5C83",
	066 => X"5947",
	067 => X"55EE",
	068 => X"5278",
	069 => X"4EE7",
	070 => X"4B3B",
	071 => X"4777",
	072 => X"439C",
	073 => X"3FAA",
	074 => X"3BA3",
	075 => X"3789",
	076 => X"335C",
	077 => X"2F1E",
	078 => X"2AD0",
	079 => X"2675",
	080 => X"220D",
	081 => X"1D99",
	082 => X"191C",
	083 => X"1497",
	084 => X"100A",
	085 => X"0B79",
	086 => X"06E3",
	087 => X"024C",
	088 => X"FDB2",
	089 => X"F91B",
	090 => X"F485",
	091 => X"EFF4",
	092 => X"EB67",
	093 => X"E6E2",
	094 => X"E265",
	095 => X"DDF1",
	096 => X"D989",
	097 => X"D52E",
	098 => X"D0E0",
	099 => X"CCA2",
	100 => X"C875",
	101 => X"C45B",
	102 => X"C054",
	103 => X"BC62",
	104 => X"B887",
	105 => X"B4C3",
	106 => X"B117",
	107 => X"AD86",
	108 => X"AA10",
	109 => X"A6B7",
	110 => X"A37B",
	111 => X"A05D",
	112 => X"9D5F",
	113 => X"9A82",
	114 => X"97C6",
	115 => X"952C",
	116 => X"92B6",
	117 => X"9063",
	118 => X"8E36",
	119 => X"8C2E",
	120 => X"8A4C",
	121 => X"8891",
	122 => X"86FE",
	123 => X"8592",
	124 => X"844F",
	125 => X"8335",
	126 => X"8244",
	127 => X"817C",
	128 => X"80DE",
	129 => X"806A",
	130 => X"8020",
	131 => X"8001",
	132 => X"800B",
	133 => X"8040",
	134 => X"809F",
	135 => X"8128",
	136 => X"81DB",
	137 => X"82B7",
	138 => X"83BD",
	139 => X"84EC",
	140 => X"8643",
	141 => X"87C3",
	142 => X"896A",
	143 => X"8B38",
	144 => X"8D2D",
	145 => X"8F48",
	146 => X"9188",
	147 => X"93EC",
	148 => X"9674",
	149 => X"991F",
	150 => X"9BEC",
	151 => X"9EDA",
	152 => X"A1E8",
	153 => X"A515",
	154 => X"A860",
	155 => X"ABC8",
	156 => X"AF4B",
	157 => X"B2EA",
	158 => X"B6A2",
	159 => X"BA71",
	160 => X"BE58",
	161 => X"C255",
	162 => X"C666",
	163 => X"CA8A",
	164 => X"CEBF",
	165 => X"D305",
	166 => X"D75A",
	167 => X"DBBC",
	168 => X"E02A",
	169 => X"E4A2",
	170 => X"E924",
	171 => X"EDAD",
	172 => X"F23C",
	173 => X"F6D0",
	174 => X"FB66",
	175 => X"0000",
	176 => X"0498",
	177 => X"092E",
	178 => X"0DC2",
	179 => X"1251",
	180 => X"16DA",
	181 => X"1B5C",
	182 => X"1FD4",
	183 => X"2442",
	184 => X"28A4",
	185 => X"2CF9",
	186 => X"313F",
	187 => X"3574",
	188 => X"3998",
	189 => X"3DA9",
	190 => X"41A6",
	191 => X"458D",
	192 => X"495C",
	193 => X"4D14",
	194 => X"50B3",
	195 => X"5436",
	196 => X"579E",
	197 => X"5AE9",
	198 => X"5E16",
	199 => X"6124",
	200 => X"6412",
	201 => X"66DF",
	202 => X"698A",
	203 => X"6C12",
	204 => X"6E76",
	205 => X"70B6",
	206 => X"72D1",
	207 => X"74C6",
	208 => X"7694",
	209 => X"783B",
	210 => X"79BB",
	211 => X"7B12",
	212 => X"7C41",
	213 => X"7D47",
	214 => X"7E23",
	215 => X"7ED6",
	216 => X"7F5F",
	217 => X"7FBE",
	218 => X"7FF3",
	219 => X"7FFD",
	220 => X"7FDE",
	221 => X"7F94",
	222 => X"7F20",
	223 => X"7E82",
	224 => X"7DBA",
	225 => X"7CC9",
	226 => X"7BAF",
	227 => X"7A6C",
	228 => X"7900",
	229 => X"776D",
	230 => X"75B2",
	231 => X"73D0",
	232 => X"71C8",
	233 => X"6F9B",
	234 => X"6D48",
	235 => X"6AD2",
	236 => X"6838",
	237 => X"657C",
	238 => X"629F",
	239 => X"5FA1",
	240 => X"5C83",
	241 => X"5947",
	242 => X"55EE",
	243 => X"5278",
	244 => X"4EE7",
	245 => X"4B3B",
	246 => X"4777",
	247 => X"439C",
	others => X"0000"
);

CONSTANT G3: hex := (
	000 => X"0000",
	001 => X"04D7",
	002 => X"09AE",
	003 => X"0E80",
	004 => X"134E",
	005 => X"1814",
	006 => X"1CD1",
	007 => X"2184",
	008 => X"262B",
	009 => X"2AC3",
	010 => X"2F4C",
	011 => X"33C3",
	012 => X"3828",
	013 => X"3C78",
	014 => X"40B2",
	015 => X"44D4",
	016 => X"48DD",
	017 => X"4CCB",
	018 => X"509D",
	019 => X"5451",
	020 => X"57E6",
	021 => X"5B5B",
	022 => X"5EAF",
	023 => X"61E0",
	024 => X"64ED",
	025 => X"67D5",
	026 => X"6A97",
	027 => X"6D32",
	028 => X"6FA5",
	029 => X"71EF",
	030 => X"740F",
	031 => X"7605",
	032 => X"77CF",
	033 => X"796D",
	034 => X"7ADF",
	035 => X"7C24",
	036 => X"7D3B",
	037 => X"7E24",
	038 => X"7EDF",
	039 => X"7F6C",
	040 => X"7FCA",
	041 => X"7FF9",
	042 => X"7FF9",
	043 => X"7FCA",
	044 => X"7F6C",
	045 => X"7EDF",
	046 => X"7E24",
	047 => X"7D3B",
	048 => X"7C24",
	049 => X"7ADF",
	050 => X"796D",
	051 => X"77CF",
	052 => X"7605",
	053 => X"740F",
	054 => X"71EF",
	055 => X"6FA5",
	056 => X"6D32",
	057 => X"6A97",
	058 => X"67D5",
	059 => X"64ED",
	060 => X"61E0",
	061 => X"5EAF",
	062 => X"5B5B",
	063 => X"57E6",
	064 => X"5451",
	065 => X"509D",
	066 => X"4CCB",
	067 => X"48DD",
	068 => X"44D4",
	069 => X"40B2",
	070 => X"3C78",
	071 => X"3828",
	072 => X"33C3",
	073 => X"2F4C",
	074 => X"2AC3",
	075 => X"262B",
	076 => X"2184",
	077 => X"1CD1",
	078 => X"1814",
	079 => X"134E",
	080 => X"0E80",
	081 => X"09AE",
	082 => X"04D7",
	083 => X"0000",
	084 => X"FB27",
	085 => X"F650",
	086 => X"F17E",
	087 => X"ECB0",
	088 => X"E7EA",
	089 => X"E32D",
	090 => X"DE7A",
	091 => X"D9D3",
	092 => X"D53B",
	093 => X"D0B2",
	094 => X"CC3B",
	095 => X"C7D6",
	096 => X"C386",
	097 => X"BF4C",
	098 => X"BB2A",
	099 => X"B721",
	100 => X"B333",
	101 => X"AF61",
	102 => X"ABAD",
	103 => X"A818",
	104 => X"A4A3",
	105 => X"A14F",
	106 => X"9E1E",
	107 => X"9B11",
	108 => X"9829",
	109 => X"9567",
	110 => X"92CC",
	111 => X"9059",
	112 => X"8E0F",
	113 => X"8BEF",
	114 => X"89F9",
	115 => X"882F",
	116 => X"8691",
	117 => X"851F",
	118 => X"83DA",
	119 => X"82C3",
	120 => X"81DA",
	121 => X"811F",
	122 => X"8092",
	123 => X"8034",
	124 => X"8005",
	125 => X"8005",
	126 => X"8034",
	127 => X"8092",
	128 => X"811F",
	129 => X"81DA",
	130 => X"82C3",
	131 => X"83DA",
	132 => X"851F",
	133 => X"8691",
	134 => X"882F",
	135 => X"89F9",
	136 => X"8BEF",
	137 => X"8E0F",
	138 => X"9059",
	139 => X"92CC",
	140 => X"9567",
	141 => X"9829",
	142 => X"9B11",
	143 => X"9E1E",
	144 => X"A14F",
	145 => X"A4A3",
	146 => X"A818",
	147 => X"ABAD",
	148 => X"AF61",
	149 => X"B333",
	150 => X"B721",
	151 => X"BB2A",
	152 => X"BF4C",
	153 => X"C386",
	154 => X"C7D6",
	155 => X"CC3B",
	156 => X"D0B2",
	157 => X"D53B",
	158 => X"D9D3",
	159 => X"DE7A",
	160 => X"E32D",
	161 => X"E7EA",
	162 => X"ECB0",
	163 => X"F17E",
	164 => X"F650",
	165 => X"FB27",
	166 => X"0000",
	167 => X"04D7",
	168 => X"09AE",
	169 => X"0E80",
	170 => X"134E",
	171 => X"1814",
	172 => X"1CD1",
	173 => X"2184",
	174 => X"262B",
	175 => X"2AC3",
	176 => X"2F4C",
	177 => X"33C3",
	178 => X"3828",
	179 => X"3C78",
	180 => X"40B2",
	181 => X"44D4",
	182 => X"48DD",
	183 => X"4CCB",
	184 => X"509D",
	185 => X"5451",
	186 => X"57E6",
	187 => X"5B5B",
	188 => X"5EAF",
	189 => X"61E0",
	190 => X"64ED",
	191 => X"67D5",
	192 => X"6A97",
	193 => X"6D32",
	194 => X"6FA5",
	195 => X"71EF",
	196 => X"740F",
	197 => X"7605",
	198 => X"77CF",
	199 => X"796D",
	200 => X"7ADF",
	201 => X"7C24",
	202 => X"7D3B",
	203 => X"7E24",
	204 => X"7EDF",
	205 => X"7F6C",
	206 => X"7FCA",
	207 => X"7FF9",
	208 => X"7FF9",
	209 => X"7FCA",
	210 => X"7F6C",
	211 => X"7EDF",
	212 => X"7E24",
	213 => X"7D3B",
	214 => X"7C24",
	215 => X"7ADF",
	216 => X"796D",
	217 => X"77CF",
	218 => X"7605",
	219 => X"740F",
	220 => X"71EF",
	221 => X"6FA5",
	222 => X"6D32",
	223 => X"6A97",
	224 => X"67D5",
	225 => X"64ED",
	226 => X"61E0",
	227 => X"5EAF",
	228 => X"5B5B",
	229 => X"57E6",
	230 => X"5451",
	231 => X"509D",
	232 => X"4CCB",
	233 => X"48DD",
	234 => X"44D4",
	235 => X"40B2",
	236 => X"3C78",
	237 => X"3828",
	238 => X"33C3",
	239 => X"2F4C",
	240 => X"2AC3",
	241 => X"262B",
	242 => X"2184",
	243 => X"1CD1",
	244 => X"1814",
	245 => X"134E",
	246 => X"0E80",
	247 => X"09AE",
	others => X"0000"
);

CONSTANT GS3: hex := (
	000 => X"0000",
	001 => X"0527",
	002 => X"0A4C",
	003 => X"0F6D",
	004 => X"1488",
	005 => X"199A",
	006 => X"1EA1",
	007 => X"239C",
	008 => X"2888",
	009 => X"2D63",
	010 => X"322B",
	011 => X"36DE",
	012 => X"3B7B",
	013 => X"3FFF",
	014 => X"4468",
	015 => X"48B5",
	016 => X"4CE4",
	017 => X"50F3",
	018 => X"54E0",
	019 => X"58AA",
	020 => X"5C4F",
	021 => X"5FCE",
	022 => X"6325",
	023 => X"6653",
	024 => X"6956",
	025 => X"6C2E",
	026 => X"6ED9",
	027 => X"7155",
	028 => X"73A3",
	029 => X"75C0",
	030 => X"77AD",
	031 => X"7968",
	032 => X"7AF1",
	033 => X"7C46",
	034 => X"7D68",
	035 => X"7E56",
	036 => X"7F10",
	037 => X"7F94",
	038 => X"7FE4",
	039 => X"7FFF",
	040 => X"7FE4",
	041 => X"7F94",
	042 => X"7F10",
	043 => X"7E56",
	044 => X"7D68",
	045 => X"7C46",
	046 => X"7AF1",
	047 => X"7968",
	048 => X"77AD",
	049 => X"75C0",
	050 => X"73A3",
	051 => X"7155",
	052 => X"6ED9",
	053 => X"6C2E",
	054 => X"6956",
	055 => X"6653",
	056 => X"6325",
	057 => X"5FCE",
	058 => X"5C4F",
	059 => X"58AA",
	060 => X"54E0",
	061 => X"50F3",
	062 => X"4CE4",
	063 => X"48B5",
	064 => X"4468",
	065 => X"3FFF",
	066 => X"3B7B",
	067 => X"36DE",
	068 => X"322B",
	069 => X"2D63",
	070 => X"2888",
	071 => X"239C",
	072 => X"1EA1",
	073 => X"199A",
	074 => X"1488",
	075 => X"0F6D",
	076 => X"0A4C",
	077 => X"0527",
	078 => X"FFFE",
	079 => X"FAD7",
	080 => X"F5B2",
	081 => X"F091",
	082 => X"EB76",
	083 => X"E664",
	084 => X"E15D",
	085 => X"DC62",
	086 => X"D776",
	087 => X"D29B",
	088 => X"CDD3",
	089 => X"C920",
	090 => X"C483",
	091 => X"BFFF",
	092 => X"BB96",
	093 => X"B749",
	094 => X"B31A",
	095 => X"AF0B",
	096 => X"AB1E",
	097 => X"A754",
	098 => X"A3AF",
	099 => X"A030",
	100 => X"9CD9",
	101 => X"99AB",
	102 => X"96A8",
	103 => X"93D0",
	104 => X"9125",
	105 => X"8EA9",
	106 => X"8C5B",
	107 => X"8A3E",
	108 => X"8851",
	109 => X"8696",
	110 => X"850D",
	111 => X"83B8",
	112 => X"8296",
	113 => X"81A8",
	114 => X"80EE",
	115 => X"806A",
	116 => X"801A",
	117 => X"8000",
	118 => X"801A",
	119 => X"806A",
	120 => X"80EE",
	121 => X"81A8",
	122 => X"8296",
	123 => X"83B8",
	124 => X"850D",
	125 => X"8696",
	126 => X"8851",
	127 => X"8A3E",
	128 => X"8C5B",
	129 => X"8EA9",
	130 => X"9125",
	131 => X"93D0",
	132 => X"96A8",
	133 => X"99AB",
	134 => X"9CD9",
	135 => X"A030",
	136 => X"A3AF",
	137 => X"A754",
	138 => X"AB1E",
	139 => X"AF0B",
	140 => X"B31A",
	141 => X"B749",
	142 => X"BB96",
	143 => X"BFFF",
	144 => X"C483",
	145 => X"C920",
	146 => X"CDD3",
	147 => X"D29B",
	148 => X"D776",
	149 => X"DC62",
	150 => X"E15D",
	151 => X"E664",
	152 => X"EB76",
	153 => X"F091",
	154 => X"F5B2",
	155 => X"FAD7",
	156 => X"0000",
	157 => X"0527",
	158 => X"0A4C",
	159 => X"0F6D",
	160 => X"1488",
	161 => X"199A",
	162 => X"1EA1",
	163 => X"239C",
	164 => X"2888",
	165 => X"2D63",
	166 => X"322B",
	167 => X"36DE",
	168 => X"3B7B",
	169 => X"3FFF",
	170 => X"4468",
	171 => X"48B5",
	172 => X"4CE4",
	173 => X"50F3",
	174 => X"54E0",
	175 => X"58AA",
	176 => X"5C4F",
	177 => X"5FCE",
	178 => X"6325",
	179 => X"6653",
	180 => X"6956",
	181 => X"6C2E",
	182 => X"6ED9",
	183 => X"7155",
	184 => X"73A3",
	185 => X"75C0",
	186 => X"77AD",
	187 => X"7968",
	188 => X"7AF1",
	189 => X"7C46",
	190 => X"7D68",
	191 => X"7E56",
	192 => X"7F10",
	193 => X"7F94",
	194 => X"7FE4",
	195 => X"7FFF",
	196 => X"7FE4",
	197 => X"7F94",
	198 => X"7F10",
	199 => X"7E56",
	200 => X"7D68",
	201 => X"7C46",
	202 => X"7AF1",
	203 => X"7968",
	204 => X"77AD",
	205 => X"75C0",
	206 => X"73A3",
	207 => X"7155",
	208 => X"6ED9",
	209 => X"6C2E",
	210 => X"6956",
	211 => X"6653",
	212 => X"6325",
	213 => X"5FCE",
	214 => X"5C4F",
	215 => X"58AA",
	216 => X"54E0",
	217 => X"50F3",
	218 => X"4CE4",
	219 => X"48B5",
	220 => X"4468",
	221 => X"3FFF",
	222 => X"3B7B",
	223 => X"36DE",
	224 => X"322B",
	225 => X"2D63",
	226 => X"2888",
	227 => X"239C",
	228 => X"1EA1",
	229 => X"199A",
	230 => X"1488",
	231 => X"0F6D",
	232 => X"0A4C",
	233 => X"0527",
	234 => X"FFFE",
	235 => X"FAD7",
	236 => X"F5B2",
	237 => X"F091",
	238 => X"EB76",
	239 => X"E664",
	240 => X"E15D",
	241 => X"DC62",
	242 => X"D776",
	243 => X"D29B",
	244 => X"CDD3",
	245 => X"C920",
	246 => X"C483",
	247 => X"BFFF",
	others => X"0000"
);

CONSTANT A3: hex := (
	000 => X"0000",
	001 => X"056E",
	002 => X"0ADA",
	003 => X"1041",
	004 => X"15A1",
	005 => X"1AF7",
	006 => X"2040",
	007 => X"257A",
	008 => X"2AA3",
	009 => X"2FB9",
	010 => X"34B8",
	011 => X"399F",
	012 => X"3E6C",
	013 => X"431B",
	014 => X"47AC",
	015 => X"4C1C",
	016 => X"5068",
	017 => X"5490",
	018 => X"5890",
	019 => X"5C68",
	020 => X"6015",
	021 => X"6395",
	022 => X"66E8",
	023 => X"6A0B",
	024 => X"6CFE",
	025 => X"6FBE",
	026 => X"724A",
	027 => X"74A2",
	028 => X"76C4",
	029 => X"78AF",
	030 => X"7A62",
	031 => X"7BDD",
	032 => X"7D1F",
	033 => X"7E27",
	034 => X"7EF5",
	035 => X"7F88",
	036 => X"7FE1",
	037 => X"7FFF",
	038 => X"7FE1",
	039 => X"7F88",
	040 => X"7EF5",
	041 => X"7E27",
	042 => X"7D1F",
	043 => X"7BDD",
	044 => X"7A62",
	045 => X"78AF",
	046 => X"76C4",
	047 => X"74A2",
	048 => X"724A",
	049 => X"6FBE",
	050 => X"6CFE",
	051 => X"6A0B",
	052 => X"66E8",
	053 => X"6395",
	054 => X"6015",
	055 => X"5C68",
	056 => X"5890",
	057 => X"5490",
	058 => X"5068",
	059 => X"4C1C",
	060 => X"47AC",
	061 => X"431B",
	062 => X"3E6C",
	063 => X"399F",
	064 => X"34B8",
	065 => X"2FB9",
	066 => X"2AA3",
	067 => X"257A",
	068 => X"2040",
	069 => X"1AF7",
	070 => X"15A1",
	071 => X"1041",
	072 => X"0ADA",
	073 => X"056E",
	074 => X"0000",
	075 => X"FA90",
	076 => X"F524",
	077 => X"EFBD",
	078 => X"EA5D",
	079 => X"E507",
	080 => X"DFBE",
	081 => X"DA84",
	082 => X"D55B",
	083 => X"D045",
	084 => X"CB46",
	085 => X"C65F",
	086 => X"C192",
	087 => X"BCE3",
	088 => X"B852",
	089 => X"B3E2",
	090 => X"AF96",
	091 => X"AB6E",
	092 => X"A76E",
	093 => X"A396",
	094 => X"9FE9",
	095 => X"9C69",
	096 => X"9916",
	097 => X"95F3",
	098 => X"9300",
	099 => X"9040",
	100 => X"8DB4",
	101 => X"8B5C",
	102 => X"893A",
	103 => X"874F",
	104 => X"859C",
	105 => X"8421",
	106 => X"82DF",
	107 => X"81D7",
	108 => X"8109",
	109 => X"8076",
	110 => X"801D",
	111 => X"8000",
	112 => X"801D",
	113 => X"8076",
	114 => X"8109",
	115 => X"81D7",
	116 => X"82DF",
	117 => X"8421",
	118 => X"859C",
	119 => X"874F",
	120 => X"893A",
	121 => X"8B5C",
	122 => X"8DB4",
	123 => X"9040",
	124 => X"9300",
	125 => X"95F3",
	126 => X"9916",
	127 => X"9C69",
	128 => X"9FE9",
	129 => X"A396",
	130 => X"A76E",
	131 => X"AB6E",
	132 => X"AF96",
	133 => X"B3E2",
	134 => X"B852",
	135 => X"BCE3",
	136 => X"C192",
	137 => X"C65F",
	138 => X"CB46",
	139 => X"D045",
	140 => X"D55B",
	141 => X"DA84",
	142 => X"DFBE",
	143 => X"E507",
	144 => X"EA5D",
	145 => X"EFBD",
	146 => X"F524",
	147 => X"FA90",
	148 => X"0000",
	149 => X"056E",
	150 => X"0ADA",
	151 => X"1041",
	152 => X"15A1",
	153 => X"1AF7",
	154 => X"2040",
	155 => X"257A",
	156 => X"2AA3",
	157 => X"2FB9",
	158 => X"34B8",
	159 => X"399F",
	160 => X"3E6C",
	161 => X"431B",
	162 => X"47AC",
	163 => X"4C1C",
	164 => X"5068",
	165 => X"5490",
	166 => X"5890",
	167 => X"5C68",
	168 => X"6015",
	169 => X"6395",
	170 => X"66E8",
	171 => X"6A0B",
	172 => X"6CFE",
	173 => X"6FBE",
	174 => X"724A",
	175 => X"74A2",
	176 => X"76C4",
	177 => X"78AF",
	178 => X"7A62",
	179 => X"7BDD",
	180 => X"7D1F",
	181 => X"7E27",
	182 => X"7EF5",
	183 => X"7F88",
	184 => X"7FE1",
	185 => X"7FFF",
	186 => X"7FE1",
	187 => X"7F88",
	188 => X"7EF5",
	189 => X"7E27",
	190 => X"7D1F",
	191 => X"7BDD",
	192 => X"7A62",
	193 => X"78AF",
	194 => X"76C4",
	195 => X"74A2",
	196 => X"724A",
	197 => X"6FBE",
	198 => X"6CFE",
	199 => X"6A0B",
	200 => X"66E8",
	201 => X"6395",
	202 => X"6015",
	203 => X"5C68",
	204 => X"5890",
	205 => X"5490",
	206 => X"5068",
	207 => X"4C1C",
	208 => X"47AC",
	209 => X"431B",
	210 => X"3E6C",
	211 => X"399F",
	212 => X"34B8",
	213 => X"2FB9",
	214 => X"2AA3",
	215 => X"257A",
	216 => X"2040",
	217 => X"1AF7",
	218 => X"15A1",
	219 => X"1041",
	220 => X"0ADA",
	221 => X"056E",
	222 => X"FFFE",
	223 => X"FA90",
	224 => X"F524",
	225 => X"EFBD",
	226 => X"EA5D",
	227 => X"E507",
	228 => X"DFBE",
	229 => X"DA84",
	230 => X"D55B",
	231 => X"D045",
	232 => X"CB46",
	233 => X"C65F",
	234 => X"C192",
	235 => X"BCE3",
	236 => X"B852",
	237 => X"B3E2",
	238 => X"AF96",
	239 => X"AB6E",
	240 => X"A76E",
	241 => X"A396",
	242 => X"9FE9",
	243 => X"9C69",
	244 => X"9916",
	245 => X"95F3",
	246 => X"9300",
	247 => X"9040",
	others => X"0000"
);

CONSTANT AS3: hex := (
	000 => X"0000",
	001 => X"05C8",
	002 => X"0B8E",
	003 => X"114D",
	004 => X"1704",
	005 => X"1CAE",
	006 => X"224A",
	007 => X"27D3",
	008 => X"2D48",
	009 => X"32A5",
	010 => X"37E8",
	011 => X"3D0D",
	012 => X"4213",
	013 => X"46F5",
	014 => X"4BB3",
	015 => X"5049",
	016 => X"54B5",
	017 => X"58F5",
	018 => X"5D07",
	019 => X"60E7",
	020 => X"6495",
	021 => X"680F",
	022 => X"6B51",
	023 => X"6E5C",
	024 => X"712D",
	025 => X"73C3",
	026 => X"761D",
	027 => X"7838",
	028 => X"7A15",
	029 => X"7BB2",
	030 => X"7D0E",
	031 => X"7E29",
	032 => X"7F02",
	033 => X"7F98",
	034 => X"7FEC",
	035 => X"7FFC",
	036 => X"7FCA",
	037 => X"7F55",
	038 => X"7E9E",
	039 => X"7DA4",
	040 => X"7C68",
	041 => X"7AEC",
	042 => X"792F",
	043 => X"7732",
	044 => X"74F8",
	045 => X"7280",
	046 => X"6FCC",
	047 => X"6CDE",
	048 => X"69B7",
	049 => X"6659",
	050 => X"62C5",
	051 => X"5EFD",
	052 => X"5B04",
	053 => X"56DB",
	054 => X"5285",
	055 => X"4E03",
	056 => X"4959",
	057 => X"4488",
	058 => X"3F94",
	059 => X"3A7E",
	060 => X"354A",
	061 => X"2FFA",
	062 => X"2A91",
	063 => X"2511",
	064 => X"1F7E",
	065 => X"19DB",
	066 => X"142A",
	067 => X"0E6F",
	068 => X"08AC",
	069 => X"02E4",
	070 => X"FD1A",
	071 => X"F752",
	072 => X"F18F",
	073 => X"EBD4",
	074 => X"E623",
	075 => X"E080",
	076 => X"DAED",
	077 => X"D56D",
	078 => X"D004",
	079 => X"CAB4",
	080 => X"C580",
	081 => X"C06A",
	082 => X"BB76",
	083 => X"B6A5",
	084 => X"B1FB",
	085 => X"AD79",
	086 => X"A923",
	087 => X"A4FA",
	088 => X"A101",
	089 => X"9D39",
	090 => X"99A5",
	091 => X"9647",
	092 => X"9320",
	093 => X"9032",
	094 => X"8D7E",
	095 => X"8B06",
	096 => X"88CC",
	097 => X"86CF",
	098 => X"8512",
	099 => X"8396",
	100 => X"825A",
	101 => X"8160",
	102 => X"80A9",
	103 => X"8034",
	104 => X"8002",
	105 => X"8012",
	106 => X"8066",
	107 => X"80FC",
	108 => X"81D5",
	109 => X"82F0",
	110 => X"844C",
	111 => X"85E9",
	112 => X"87C6",
	113 => X"89E1",
	114 => X"8C3B",
	115 => X"8ED1",
	116 => X"91A2",
	117 => X"94AD",
	118 => X"97EF",
	119 => X"9B69",
	120 => X"9F17",
	121 => X"A2F7",
	122 => X"A709",
	123 => X"AB49",
	124 => X"AFB5",
	125 => X"B44B",
	126 => X"B909",
	127 => X"BDEB",
	128 => X"C2F1",
	129 => X"C816",
	130 => X"CD59",
	131 => X"D2B6",
	132 => X"D82B",
	133 => X"DDB4",
	134 => X"E350",
	135 => X"E8FA",
	136 => X"EEB1",
	137 => X"F470",
	138 => X"FA36",
	139 => X"FFFE",
	140 => X"05C8",
	141 => X"0B8E",
	142 => X"114D",
	143 => X"1704",
	144 => X"1CAE",
	145 => X"224A",
	146 => X"27D3",
	147 => X"2D48",
	148 => X"32A5",
	149 => X"37E8",
	150 => X"3D0D",
	151 => X"4213",
	152 => X"46F5",
	153 => X"4BB3",
	154 => X"5049",
	155 => X"54B5",
	156 => X"58F5",
	157 => X"5D07",
	158 => X"60E7",
	159 => X"6495",
	160 => X"680F",
	161 => X"6B51",
	162 => X"6E5C",
	163 => X"712D",
	164 => X"73C3",
	165 => X"761D",
	166 => X"7838",
	167 => X"7A15",
	168 => X"7BB2",
	169 => X"7D0E",
	170 => X"7E29",
	171 => X"7F02",
	172 => X"7F98",
	173 => X"7FEC",
	174 => X"7FFC",
	175 => X"7FCA",
	176 => X"7F55",
	177 => X"7E9E",
	178 => X"7DA4",
	179 => X"7C68",
	180 => X"7AEC",
	181 => X"792F",
	182 => X"7732",
	183 => X"74F8",
	184 => X"7280",
	185 => X"6FCC",
	186 => X"6CDE",
	187 => X"69B7",
	188 => X"6659",
	189 => X"62C5",
	190 => X"5EFD",
	191 => X"5B04",
	192 => X"56DB",
	193 => X"5285",
	194 => X"4E03",
	195 => X"4959",
	196 => X"4488",
	197 => X"3F94",
	198 => X"3A7E",
	199 => X"354A",
	200 => X"2FFA",
	201 => X"2A91",
	202 => X"2511",
	203 => X"1F7E",
	204 => X"19DB",
	205 => X"142A",
	206 => X"0E6F",
	207 => X"08AC",
	208 => X"02E4",
	209 => X"FD1A",
	210 => X"F752",
	211 => X"F18F",
	212 => X"EBD4",
	213 => X"E623",
	214 => X"E080",
	215 => X"DAED",
	216 => X"D56D",
	217 => X"D004",
	218 => X"CAB4",
	219 => X"C580",
	220 => X"C06A",
	221 => X"BB76",
	222 => X"B6A5",
	223 => X"B1FB",
	224 => X"AD79",
	225 => X"A923",
	226 => X"A4FA",
	227 => X"A101",
	228 => X"9D39",
	229 => X"99A5",
	230 => X"9647",
	231 => X"9320",
	232 => X"9032",
	233 => X"8D7E",
	234 => X"8B06",
	235 => X"88CC",
	236 => X"86CF",
	237 => X"8512",
	238 => X"8396",
	239 => X"825A",
	240 => X"8160",
	241 => X"80A9",
	242 => X"8034",
	243 => X"8002",
	244 => X"8012",
	245 => X"8066",
	246 => X"80FC",
	247 => X"81D5",
	others => X"0000"
);

CONSTANT B3: hex := (
	000 => X"0000",
	001 => X"0623",
	002 => X"0C42",
	003 => X"125A",
	004 => X"1867",
	005 => X"1E66",
	006 => X"2454",
	007 => X"2A2B",
	008 => X"2FEA",
	009 => X"358D",
	010 => X"3B10",
	011 => X"4070",
	012 => X"45AB",
	013 => X"4ABC",
	014 => X"4FA1",
	015 => X"5458",
	016 => X"58DD",
	017 => X"5D2D",
	018 => X"6147",
	019 => X"6527",
	020 => X"68CC",
	021 => X"6C33",
	022 => X"6F5B",
	023 => X"7240",
	024 => X"74E3",
	025 => X"7741",
	026 => X"7958",
	027 => X"7B28",
	028 => X"7CB0",
	029 => X"7DEE",
	030 => X"7EE2",
	031 => X"7F8B",
	032 => X"7FE9",
	033 => X"7FFC",
	034 => X"7FC4",
	035 => X"7F40",
	036 => X"7E71",
	037 => X"7D58",
	038 => X"7BF5",
	039 => X"7A49",
	040 => X"7855",
	041 => X"761B",
	042 => X"739A",
	043 => X"70D6",
	044 => X"6DCF",
	045 => X"6A88",
	046 => X"6701",
	047 => X"633E",
	048 => X"5F41",
	049 => X"5B0C",
	050 => X"56A1",
	051 => X"5203",
	052 => X"4D34",
	053 => X"4839",
	054 => X"4312",
	055 => X"3DC5",
	056 => X"3853",
	057 => X"32BF",
	058 => X"2D0E",
	059 => X"2742",
	060 => X"215F",
	061 => X"1B69",
	062 => X"1562",
	063 => X"0F4F",
	064 => X"0933",
	065 => X"0311",
	066 => X"FCED",
	067 => X"F6CB",
	068 => X"F0AF",
	069 => X"EA9C",
	070 => X"E495",
	071 => X"DE9F",
	072 => X"D8BC",
	073 => X"D2F0",
	074 => X"CD3F",
	075 => X"C7AB",
	076 => X"C239",
	077 => X"BCEC",
	078 => X"B7C5",
	079 => X"B2CA",
	080 => X"ADFB",
	081 => X"A95D",
	082 => X"A4F2",
	083 => X"A0BD",
	084 => X"9CC0",
	085 => X"98FD",
	086 => X"9576",
	087 => X"922F",
	088 => X"8F28",
	089 => X"8C64",
	090 => X"89E3",
	091 => X"87A9",
	092 => X"85B5",
	093 => X"8409",
	094 => X"82A6",
	095 => X"818D",
	096 => X"80BE",
	097 => X"803A",
	098 => X"8002",
	099 => X"8015",
	100 => X"8073",
	101 => X"811C",
	102 => X"8210",
	103 => X"834E",
	104 => X"84D6",
	105 => X"86A6",
	106 => X"88BD",
	107 => X"8B1B",
	108 => X"8DBE",
	109 => X"90A3",
	110 => X"93CB",
	111 => X"9732",
	112 => X"9AD7",
	113 => X"9EB7",
	114 => X"A2D1",
	115 => X"A721",
	116 => X"ABA6",
	117 => X"B05D",
	118 => X"B542",
	119 => X"BA53",
	120 => X"BF8E",
	121 => X"C4EE",
	122 => X"CA71",
	123 => X"D014",
	124 => X"D5D3",
	125 => X"DBAA",
	126 => X"E198",
	127 => X"E797",
	128 => X"EDA4",
	129 => X"F3BC",
	130 => X"F9DB",
	131 => X"FFFE",
	132 => X"0623",
	133 => X"0C42",
	134 => X"125A",
	135 => X"1867",
	136 => X"1E66",
	137 => X"2454",
	138 => X"2A2B",
	139 => X"2FEA",
	140 => X"358D",
	141 => X"3B10",
	142 => X"4070",
	143 => X"45AB",
	144 => X"4ABC",
	145 => X"4FA1",
	146 => X"5458",
	147 => X"58DD",
	148 => X"5D2D",
	149 => X"6147",
	150 => X"6527",
	151 => X"68CC",
	152 => X"6C33",
	153 => X"6F5B",
	154 => X"7240",
	155 => X"74E3",
	156 => X"7741",
	157 => X"7958",
	158 => X"7B28",
	159 => X"7CB0",
	160 => X"7DEE",
	161 => X"7EE2",
	162 => X"7F8B",
	163 => X"7FE9",
	164 => X"7FFC",
	165 => X"7FC4",
	166 => X"7F40",
	167 => X"7E71",
	168 => X"7D58",
	169 => X"7BF5",
	170 => X"7A49",
	171 => X"7855",
	172 => X"761B",
	173 => X"739A",
	174 => X"70D6",
	175 => X"6DCF",
	176 => X"6A88",
	177 => X"6701",
	178 => X"633E",
	179 => X"5F41",
	180 => X"5B0C",
	181 => X"56A1",
	182 => X"5203",
	183 => X"4D34",
	184 => X"4839",
	185 => X"4312",
	186 => X"3DC5",
	187 => X"3853",
	188 => X"32BF",
	189 => X"2D0E",
	190 => X"2742",
	191 => X"215F",
	192 => X"1B69",
	193 => X"1562",
	194 => X"0F4F",
	195 => X"0933",
	196 => X"0311",
	197 => X"FCED",
	198 => X"F6CB",
	199 => X"F0AF",
	200 => X"EA9C",
	201 => X"E495",
	202 => X"DE9F",
	203 => X"D8BC",
	204 => X"D2F0",
	205 => X"CD3F",
	206 => X"C7AB",
	207 => X"C239",
	208 => X"BCEC",
	209 => X"B7C5",
	210 => X"B2CA",
	211 => X"ADFB",
	212 => X"A95D",
	213 => X"A4F2",
	214 => X"A0BD",
	215 => X"9CC0",
	216 => X"98FD",
	217 => X"9576",
	218 => X"922F",
	219 => X"8F28",
	220 => X"8C64",
	221 => X"89E3",
	222 => X"87A9",
	223 => X"85B5",
	224 => X"8409",
	225 => X"82A6",
	226 => X"818D",
	227 => X"80BE",
	228 => X"803A",
	229 => X"8002",
	230 => X"8015",
	231 => X"8073",
	232 => X"811C",
	233 => X"8210",
	234 => X"834E",
	235 => X"84D6",
	236 => X"86A6",
	237 => X"88BD",
	238 => X"8B1B",
	239 => X"8DBE",
	240 => X"90A3",
	241 => X"93CB",
	242 => X"9732",
	243 => X"9AD7",
	244 => X"9EB7",
	245 => X"A2D1",
	246 => X"A721",
	247 => X"ABA6",
	others => X"0000"
);

CONSTANT C4: hex := (
	000 => X"0000",
	001 => X"067B",
	002 => X"0CF2",
	003 => X"1361",
	004 => X"19C3",
	005 => X"2015",
	006 => X"2651",
	007 => X"2C74",
	008 => X"3279",
	009 => X"385E",
	010 => X"3E1D",
	011 => X"43B4",
	012 => X"491E",
	013 => X"4E58",
	014 => X"535F",
	015 => X"582F",
	016 => X"5CC5",
	017 => X"611E",
	018 => X"6537",
	019 => X"690D",
	020 => X"6C9F",
	021 => X"6FE9",
	022 => X"72EA",
	023 => X"759F",
	024 => X"7807",
	025 => X"7A20",
	026 => X"7BE8",
	027 => X"7D60",
	028 => X"7E85",
	029 => X"7F56",
	030 => X"7FD4",
	031 => X"7FFF",
	032 => X"7FD4",
	033 => X"7F56",
	034 => X"7E85",
	035 => X"7D60",
	036 => X"7BE8",
	037 => X"7A20",
	038 => X"7807",
	039 => X"759F",
	040 => X"72EA",
	041 => X"6FE9",
	042 => X"6C9F",
	043 => X"690D",
	044 => X"6537",
	045 => X"611E",
	046 => X"5CC5",
	047 => X"582F",
	048 => X"535F",
	049 => X"4E58",
	050 => X"491E",
	051 => X"43B4",
	052 => X"3E1D",
	053 => X"385E",
	054 => X"3279",
	055 => X"2C74",
	056 => X"2651",
	057 => X"2015",
	058 => X"19C3",
	059 => X"1361",
	060 => X"0CF2",
	061 => X"067B",
	062 => X"FFFE",
	063 => X"F983",
	064 => X"F30C",
	065 => X"EC9D",
	066 => X"E63B",
	067 => X"DFE9",
	068 => X"D9AD",
	069 => X"D38A",
	070 => X"CD85",
	071 => X"C7A0",
	072 => X"C1E1",
	073 => X"BC4A",
	074 => X"B6E0",
	075 => X"B1A6",
	076 => X"AC9F",
	077 => X"A7CF",
	078 => X"A339",
	079 => X"9EE0",
	080 => X"9AC7",
	081 => X"96F1",
	082 => X"935F",
	083 => X"9015",
	084 => X"8D14",
	085 => X"8A5F",
	086 => X"87F7",
	087 => X"85DE",
	088 => X"8416",
	089 => X"829E",
	090 => X"8179",
	091 => X"80A8",
	092 => X"802A",
	093 => X"8000",
	094 => X"802A",
	095 => X"80A8",
	096 => X"8179",
	097 => X"829E",
	098 => X"8416",
	099 => X"85DE",
	100 => X"87F7",
	101 => X"8A5F",
	102 => X"8D14",
	103 => X"9015",
	104 => X"935F",
	105 => X"96F1",
	106 => X"9AC7",
	107 => X"9EE0",
	108 => X"A339",
	109 => X"A7CF",
	110 => X"AC9F",
	111 => X"B1A6",
	112 => X"B6E0",
	113 => X"BC4A",
	114 => X"C1E1",
	115 => X"C7A0",
	116 => X"CD85",
	117 => X"D38A",
	118 => X"D9AD",
	119 => X"DFE9",
	120 => X"E63B",
	121 => X"EC9D",
	122 => X"F30C",
	123 => X"F983",
	124 => X"FFFE",
	125 => X"067B",
	126 => X"0CF2",
	127 => X"1361",
	128 => X"19C3",
	129 => X"2015",
	130 => X"2651",
	131 => X"2C74",
	132 => X"3279",
	133 => X"385E",
	134 => X"3E1D",
	135 => X"43B4",
	136 => X"491E",
	137 => X"4E58",
	138 => X"535F",
	139 => X"582F",
	140 => X"5CC5",
	141 => X"611E",
	142 => X"6537",
	143 => X"690D",
	144 => X"6C9F",
	145 => X"6FE9",
	146 => X"72EA",
	147 => X"759F",
	148 => X"7807",
	149 => X"7A20",
	150 => X"7BE8",
	151 => X"7D60",
	152 => X"7E85",
	153 => X"7F56",
	154 => X"7FD4",
	155 => X"7FFF",
	156 => X"7FD4",
	157 => X"7F56",
	158 => X"7E85",
	159 => X"7D60",
	160 => X"7BE8",
	161 => X"7A20",
	162 => X"7807",
	163 => X"759F",
	164 => X"72EA",
	165 => X"6FE9",
	166 => X"6C9F",
	167 => X"690D",
	168 => X"6537",
	169 => X"611E",
	170 => X"5CC5",
	171 => X"582F",
	172 => X"535F",
	173 => X"4E58",
	174 => X"491E",
	175 => X"43B4",
	176 => X"3E1D",
	177 => X"385E",
	178 => X"3279",
	179 => X"2C74",
	180 => X"2651",
	181 => X"2015",
	182 => X"19C3",
	183 => X"1361",
	184 => X"0CF2",
	185 => X"067B",
	186 => X"0000",
	187 => X"F983",
	188 => X"F30C",
	189 => X"EC9D",
	190 => X"E63B",
	191 => X"DFE9",
	192 => X"D9AD",
	193 => X"D38A",
	194 => X"CD85",
	195 => X"C7A0",
	196 => X"C1E1",
	197 => X"BC4A",
	198 => X"B6E0",
	199 => X"B1A6",
	200 => X"AC9F",
	201 => X"A7CF",
	202 => X"A339",
	203 => X"9EE0",
	204 => X"9AC7",
	205 => X"96F1",
	206 => X"935F",
	207 => X"9015",
	208 => X"8D14",
	209 => X"8A5F",
	210 => X"87F7",
	211 => X"85DE",
	212 => X"8416",
	213 => X"829E",
	214 => X"8179",
	215 => X"80A8",
	216 => X"802A",
	217 => X"8000",
	218 => X"802A",
	219 => X"80A8",
	220 => X"8179",
	221 => X"829E",
	222 => X"8416",
	223 => X"85DE",
	224 => X"87F7",
	225 => X"8A5F",
	226 => X"8D14",
	227 => X"9015",
	228 => X"935F",
	229 => X"96F1",
	230 => X"9AC7",
	231 => X"9EE0",
	232 => X"A339",
	233 => X"A7CF",
	234 => X"AC9F",
	235 => X"B1A6",
	236 => X"B6E0",
	237 => X"BC4A",
	238 => X"C1E1",
	239 => X"C7A0",
	240 => X"CD85",
	241 => X"D38A",
	242 => X"D9AD",
	243 => X"DFE9",
	244 => X"E63B",
	245 => X"EC9D",
	246 => X"F30C",
	247 => X"F983",
	others => X"0000"
);

CONSTANT CS4: hex := (
	000 => X"0000",
	001 => X"06DE",
	002 => X"0DB8",
	003 => X"1488",
	004 => X"1B48",
	005 => X"21F4",
	006 => X"2888",
	007 => X"2EFD",
	008 => X"3550",
	009 => X"3B7B",
	010 => X"417A",
	011 => X"474A",
	012 => X"4CE4",
	013 => X"5246",
	014 => X"576B",
	015 => X"5C4F",
	016 => X"60EF",
	017 => X"6548",
	018 => X"6956",
	019 => X"6D16",
	020 => X"7086",
	021 => X"73A3",
	022 => X"766A",
	023 => X"78DA",
	024 => X"7AF1",
	025 => X"7CAD",
	026 => X"7E0D",
	027 => X"7F10",
	028 => X"7FB5",
	029 => X"7FFC",
	030 => X"7FE4",
	031 => X"7F6E",
	032 => X"7E9A",
	033 => X"7D68",
	034 => X"7BDA",
	035 => X"79F1",
	036 => X"77AD",
	037 => X"7511",
	038 => X"721F",
	039 => X"6ED9",
	040 => X"6B40",
	041 => X"6759",
	042 => X"6325",
	043 => X"5EA8",
	044 => X"59E5",
	045 => X"54E0",
	046 => X"4F9C",
	047 => X"4A1E",
	048 => X"4468",
	049 => X"3E81",
	050 => X"386B",
	051 => X"322B",
	052 => X"2BC6",
	053 => X"2542",
	054 => X"1EA1",
	055 => X"17EA",
	056 => X"1121",
	057 => X"0A4C",
	058 => X"036F",
	059 => X"FC8F",
	060 => X"F5B2",
	061 => X"EEDD",
	062 => X"E814",
	063 => X"E15D",
	064 => X"DABC",
	065 => X"D438",
	066 => X"CDD3",
	067 => X"C793",
	068 => X"C17D",
	069 => X"BB96",
	070 => X"B5E0",
	071 => X"B062",
	072 => X"AB1E",
	073 => X"A619",
	074 => X"A156",
	075 => X"9CD9",
	076 => X"98A5",
	077 => X"94BE",
	078 => X"9125",
	079 => X"8DDF",
	080 => X"8AED",
	081 => X"8851",
	082 => X"860D",
	083 => X"8424",
	084 => X"8296",
	085 => X"8164",
	086 => X"8090",
	087 => X"801A",
	088 => X"8002",
	089 => X"8049",
	090 => X"80EE",
	091 => X"81F1",
	092 => X"8351",
	093 => X"850D",
	094 => X"8724",
	095 => X"8994",
	096 => X"8C5B",
	097 => X"8F78",
	098 => X"92E8",
	099 => X"96A8",
	100 => X"9AB6",
	101 => X"9F0F",
	102 => X"A3AF",
	103 => X"A893",
	104 => X"ADB8",
	105 => X"B31A",
	106 => X"B8B4",
	107 => X"BE84",
	108 => X"C483",
	109 => X"CAAE",
	110 => X"D101",
	111 => X"D776",
	112 => X"DE0A",
	113 => X"E4B6",
	114 => X"EB76",
	115 => X"F246",
	116 => X"F920",
	117 => X"0000",
	118 => X"06DE",
	119 => X"0DB8",
	120 => X"1488",
	121 => X"1B48",
	122 => X"21F4",
	123 => X"2888",
	124 => X"2EFD",
	125 => X"3550",
	126 => X"3B7B",
	127 => X"417A",
	128 => X"474A",
	129 => X"4CE4",
	130 => X"5246",
	131 => X"576B",
	132 => X"5C4F",
	133 => X"60EF",
	134 => X"6548",
	135 => X"6956",
	136 => X"6D16",
	137 => X"7086",
	138 => X"73A3",
	139 => X"766A",
	140 => X"78DA",
	141 => X"7AF1",
	142 => X"7CAD",
	143 => X"7E0D",
	144 => X"7F10",
	145 => X"7FB5",
	146 => X"7FFC",
	147 => X"7FE4",
	148 => X"7F6E",
	149 => X"7E9A",
	150 => X"7D68",
	151 => X"7BDA",
	152 => X"79F1",
	153 => X"77AD",
	154 => X"7511",
	155 => X"721F",
	156 => X"6ED9",
	157 => X"6B40",
	158 => X"6759",
	159 => X"6325",
	160 => X"5EA8",
	161 => X"59E5",
	162 => X"54E0",
	163 => X"4F9C",
	164 => X"4A1E",
	165 => X"4468",
	166 => X"3E81",
	167 => X"386B",
	168 => X"322B",
	169 => X"2BC6",
	170 => X"2542",
	171 => X"1EA1",
	172 => X"17EA",
	173 => X"1121",
	174 => X"0A4C",
	175 => X"036F",
	176 => X"FC8F",
	177 => X"F5B2",
	178 => X"EEDD",
	179 => X"E814",
	180 => X"E15D",
	181 => X"DABC",
	182 => X"D438",
	183 => X"CDD3",
	184 => X"C793",
	185 => X"C17D",
	186 => X"BB96",
	187 => X"B5E0",
	188 => X"B062",
	189 => X"AB1E",
	190 => X"A619",
	191 => X"A156",
	192 => X"9CD9",
	193 => X"98A5",
	194 => X"94BE",
	195 => X"9125",
	196 => X"8DDF",
	197 => X"8AED",
	198 => X"8851",
	199 => X"860D",
	200 => X"8424",
	201 => X"8296",
	202 => X"8164",
	203 => X"8090",
	204 => X"801A",
	205 => X"8002",
	206 => X"8049",
	207 => X"80EE",
	208 => X"81F1",
	209 => X"8351",
	210 => X"850D",
	211 => X"8724",
	212 => X"8994",
	213 => X"8C5B",
	214 => X"8F78",
	215 => X"92E8",
	216 => X"96A8",
	217 => X"9AB6",
	218 => X"9F0F",
	219 => X"A3AF",
	220 => X"A893",
	221 => X"ADB8",
	222 => X"B31A",
	223 => X"B8B4",
	224 => X"BE84",
	225 => X"C483",
	226 => X"CAAE",
	227 => X"D101",
	228 => X"D776",
	229 => X"DE0A",
	230 => X"E4B6",
	231 => X"EB76",
	232 => X"F246",
	233 => X"F920",
	234 => X"0000",
	235 => X"06DE",
	236 => X"0DB8",
	237 => X"1488",
	238 => X"1B48",
	239 => X"21F4",
	240 => X"2888",
	241 => X"2EFD",
	242 => X"3550",
	243 => X"3B7B",
	244 => X"417A",
	245 => X"474A",
	246 => X"4CE4",
	247 => X"5246",
	others => X"0000"
);

CONSTANT D4: hex := (
	000 => X"0000",
	001 => X"074E",
	002 => X"0E97",
	003 => X"15D3",
	004 => X"1CFD",
	005 => X"240F",
	006 => X"2B03",
	007 => X"31D3",
	008 => X"3879",
	009 => X"3EF0",
	010 => X"4533",
	011 => X"4B3B",
	012 => X"5105",
	013 => X"568C",
	014 => X"5BCA",
	015 => X"60BB",
	016 => X"655C",
	017 => X"69A8",
	018 => X"6D9B",
	019 => X"7134",
	020 => X"746D",
	021 => X"7746",
	022 => X"79BB",
	023 => X"7BCA",
	024 => X"7D72",
	025 => X"7EB1",
	026 => X"7F86",
	027 => X"7FF1",
	028 => X"7FF1",
	029 => X"7F86",
	030 => X"7EB1",
	031 => X"7D72",
	032 => X"7BCA",
	033 => X"79BB",
	034 => X"7746",
	035 => X"746D",
	036 => X"7134",
	037 => X"6D9B",
	038 => X"69A8",
	039 => X"655C",
	040 => X"60BB",
	041 => X"5BCA",
	042 => X"568C",
	043 => X"5105",
	044 => X"4B3B",
	045 => X"4533",
	046 => X"3EF0",
	047 => X"3879",
	048 => X"31D3",
	049 => X"2B03",
	050 => X"240F",
	051 => X"1CFD",
	052 => X"15D3",
	053 => X"0E97",
	054 => X"074E",
	055 => X"0000",
	056 => X"F8B0",
	057 => X"F167",
	058 => X"EA2B",
	059 => X"E301",
	060 => X"DBEF",
	061 => X"D4FB",
	062 => X"CE2B",
	063 => X"C785",
	064 => X"C10E",
	065 => X"BACB",
	066 => X"B4C3",
	067 => X"AEF9",
	068 => X"A972",
	069 => X"A434",
	070 => X"9F43",
	071 => X"9AA2",
	072 => X"9656",
	073 => X"9263",
	074 => X"8ECA",
	075 => X"8B91",
	076 => X"88B8",
	077 => X"8643",
	078 => X"8434",
	079 => X"828C",
	080 => X"814D",
	081 => X"8078",
	082 => X"800D",
	083 => X"800D",
	084 => X"8078",
	085 => X"814D",
	086 => X"828C",
	087 => X"8434",
	088 => X"8643",
	089 => X"88B8",
	090 => X"8B91",
	091 => X"8ECA",
	092 => X"9263",
	093 => X"9656",
	094 => X"9AA2",
	095 => X"9F43",
	096 => X"A434",
	097 => X"A972",
	098 => X"AEF9",
	099 => X"B4C3",
	100 => X"BACB",
	101 => X"C10E",
	102 => X"C785",
	103 => X"CE2B",
	104 => X"D4FB",
	105 => X"DBEF",
	106 => X"E301",
	107 => X"EA2B",
	108 => X"F167",
	109 => X"F8B0",
	110 => X"FFFE",
	111 => X"074E",
	112 => X"0E97",
	113 => X"15D3",
	114 => X"1CFD",
	115 => X"240F",
	116 => X"2B03",
	117 => X"31D3",
	118 => X"3879",
	119 => X"3EF0",
	120 => X"4533",
	121 => X"4B3B",
	122 => X"5105",
	123 => X"568C",
	124 => X"5BCA",
	125 => X"60BB",
	126 => X"655C",
	127 => X"69A8",
	128 => X"6D9B",
	129 => X"7134",
	130 => X"746D",
	131 => X"7746",
	132 => X"79BB",
	133 => X"7BCA",
	134 => X"7D72",
	135 => X"7EB1",
	136 => X"7F86",
	137 => X"7FF1",
	138 => X"7FF1",
	139 => X"7F86",
	140 => X"7EB1",
	141 => X"7D72",
	142 => X"7BCA",
	143 => X"79BB",
	144 => X"7746",
	145 => X"746D",
	146 => X"7134",
	147 => X"6D9B",
	148 => X"69A8",
	149 => X"655C",
	150 => X"60BB",
	151 => X"5BCA",
	152 => X"568C",
	153 => X"5105",
	154 => X"4B3B",
	155 => X"4533",
	156 => X"3EF0",
	157 => X"3879",
	158 => X"31D3",
	159 => X"2B03",
	160 => X"240F",
	161 => X"1CFD",
	162 => X"15D3",
	163 => X"0E97",
	164 => X"074E",
	165 => X"0000",
	166 => X"F8B0",
	167 => X"F167",
	168 => X"EA2B",
	169 => X"E301",
	170 => X"DBEF",
	171 => X"D4FB",
	172 => X"CE2B",
	173 => X"C785",
	174 => X"C10E",
	175 => X"BACB",
	176 => X"B4C3",
	177 => X"AEF9",
	178 => X"A972",
	179 => X"A434",
	180 => X"9F43",
	181 => X"9AA2",
	182 => X"9656",
	183 => X"9263",
	184 => X"8ECA",
	185 => X"8B91",
	186 => X"88B8",
	187 => X"8643",
	188 => X"8434",
	189 => X"828C",
	190 => X"814D",
	191 => X"8078",
	192 => X"800D",
	193 => X"800D",
	194 => X"8078",
	195 => X"814D",
	196 => X"828C",
	197 => X"8434",
	198 => X"8643",
	199 => X"88B8",
	200 => X"8B91",
	201 => X"8ECA",
	202 => X"9263",
	203 => X"9656",
	204 => X"9AA2",
	205 => X"9F43",
	206 => X"A434",
	207 => X"A972",
	208 => X"AEF9",
	209 => X"B4C3",
	210 => X"BACB",
	211 => X"C10E",
	212 => X"C785",
	213 => X"CE2B",
	214 => X"D4FB",
	215 => X"DBEF",
	216 => X"E301",
	217 => X"EA2B",
	218 => X"F167",
	219 => X"F8B0",
	220 => X"FFFE",
	221 => X"074E",
	222 => X"0E97",
	223 => X"15D3",
	224 => X"1CFD",
	225 => X"240F",
	226 => X"2B03",
	227 => X"31D3",
	228 => X"3879",
	229 => X"3EF0",
	230 => X"4533",
	231 => X"4B3B",
	232 => X"5105",
	233 => X"568C",
	234 => X"5BCA",
	235 => X"60BB",
	236 => X"655C",
	237 => X"69A8",
	238 => X"6D9B",
	239 => X"7134",
	240 => X"746D",
	241 => X"7746",
	242 => X"79BB",
	243 => X"7BCA",
	244 => X"7D72",
	245 => X"7EB1",
	246 => X"7F86",
	247 => X"7FF1",
	others => X"0000"
);

CONSTANT DS4: hex := (
	000 => X"0000",
	001 => X"07BA",
	002 => X"0F6D",
	003 => X"1712",
	004 => X"1EA1",
	005 => X"2614",
	006 => X"2D63",
	007 => X"3487",
	008 => X"3B7B",
	009 => X"4237",
	010 => X"48B5",
	011 => X"4EF0",
	012 => X"54E0",
	013 => X"5A81",
	014 => X"5FCE",
	015 => X"64C1",
	016 => X"6956",
	017 => X"6D89",
	018 => X"7155",
	019 => X"74B8",
	020 => X"77AD",
	021 => X"7A33",
	022 => X"7C46",
	023 => X"7DE6",
	024 => X"7F10",
	025 => X"7FC3",
	026 => X"7FFF",
	027 => X"7FC3",
	028 => X"7F10",
	029 => X"7DE6",
	030 => X"7C46",
	031 => X"7A33",
	032 => X"77AD",
	033 => X"74B8",
	034 => X"7155",
	035 => X"6D89",
	036 => X"6956",
	037 => X"64C1",
	038 => X"5FCE",
	039 => X"5A81",
	040 => X"54E0",
	041 => X"4EF0",
	042 => X"48B5",
	043 => X"4237",
	044 => X"3B7B",
	045 => X"3487",
	046 => X"2D63",
	047 => X"2614",
	048 => X"1EA1",
	049 => X"1712",
	050 => X"0F6D",
	051 => X"07BA",
	052 => X"0000",
	053 => X"F844",
	054 => X"F091",
	055 => X"E8EC",
	056 => X"E15D",
	057 => X"D9EA",
	058 => X"D29B",
	059 => X"CB77",
	060 => X"C483",
	061 => X"BDC7",
	062 => X"B749",
	063 => X"B10E",
	064 => X"AB1E",
	065 => X"A57D",
	066 => X"A030",
	067 => X"9B3D",
	068 => X"96A8",
	069 => X"9275",
	070 => X"8EA9",
	071 => X"8B46",
	072 => X"8851",
	073 => X"85CB",
	074 => X"83B8",
	075 => X"8218",
	076 => X"80EE",
	077 => X"803B",
	078 => X"8000",
	079 => X"803B",
	080 => X"80EE",
	081 => X"8218",
	082 => X"83B8",
	083 => X"85CB",
	084 => X"8851",
	085 => X"8B46",
	086 => X"8EA9",
	087 => X"9275",
	088 => X"96A8",
	089 => X"9B3D",
	090 => X"A030",
	091 => X"A57D",
	092 => X"AB1E",
	093 => X"B10E",
	094 => X"B749",
	095 => X"BDC7",
	096 => X"C483",
	097 => X"CB77",
	098 => X"D29B",
	099 => X"D9EA",
	100 => X"E15D",
	101 => X"E8EC",
	102 => X"F091",
	103 => X"F844",
	104 => X"FFFE",
	105 => X"07BA",
	106 => X"0F6D",
	107 => X"1712",
	108 => X"1EA1",
	109 => X"2614",
	110 => X"2D63",
	111 => X"3487",
	112 => X"3B7B",
	113 => X"4237",
	114 => X"48B5",
	115 => X"4EF0",
	116 => X"54E0",
	117 => X"5A81",
	118 => X"5FCE",
	119 => X"64C1",
	120 => X"6956",
	121 => X"6D89",
	122 => X"7155",
	123 => X"74B8",
	124 => X"77AD",
	125 => X"7A33",
	126 => X"7C46",
	127 => X"7DE6",
	128 => X"7F10",
	129 => X"7FC3",
	130 => X"7FFF",
	131 => X"7FC3",
	132 => X"7F10",
	133 => X"7DE6",
	134 => X"7C46",
	135 => X"7A33",
	136 => X"77AD",
	137 => X"74B8",
	138 => X"7155",
	139 => X"6D89",
	140 => X"6956",
	141 => X"64C1",
	142 => X"5FCE",
	143 => X"5A81",
	144 => X"54E0",
	145 => X"4EF0",
	146 => X"48B5",
	147 => X"4237",
	148 => X"3B7B",
	149 => X"3487",
	150 => X"2D63",
	151 => X"2614",
	152 => X"1EA1",
	153 => X"1712",
	154 => X"0F6D",
	155 => X"07BA",
	156 => X"0000",
	157 => X"F844",
	158 => X"F091",
	159 => X"E8EC",
	160 => X"E15D",
	161 => X"D9EA",
	162 => X"D29B",
	163 => X"CB77",
	164 => X"C483",
	165 => X"BDC7",
	166 => X"B749",
	167 => X"B10E",
	168 => X"AB1E",
	169 => X"A57D",
	170 => X"A030",
	171 => X"9B3D",
	172 => X"96A8",
	173 => X"9275",
	174 => X"8EA9",
	175 => X"8B46",
	176 => X"8851",
	177 => X"85CB",
	178 => X"83B8",
	179 => X"8218",
	180 => X"80EE",
	181 => X"803B",
	182 => X"8000",
	183 => X"803B",
	184 => X"80EE",
	185 => X"8218",
	186 => X"83B8",
	187 => X"85CB",
	188 => X"8851",
	189 => X"8B46",
	190 => X"8EA9",
	191 => X"9275",
	192 => X"96A8",
	193 => X"9B3D",
	194 => X"A030",
	195 => X"A57D",
	196 => X"AB1E",
	197 => X"B10E",
	198 => X"B749",
	199 => X"BDC7",
	200 => X"C483",
	201 => X"CB77",
	202 => X"D29B",
	203 => X"D9EA",
	204 => X"E15D",
	205 => X"E8EC",
	206 => X"F091",
	207 => X"F844",
	208 => X"FFFE",
	209 => X"07BA",
	210 => X"0F6D",
	211 => X"1712",
	212 => X"1EA1",
	213 => X"2614",
	214 => X"2D63",
	215 => X"3487",
	216 => X"3B7B",
	217 => X"4237",
	218 => X"48B5",
	219 => X"4EF0",
	220 => X"54E0",
	221 => X"5A81",
	222 => X"5FCE",
	223 => X"64C1",
	224 => X"6956",
	225 => X"6D89",
	226 => X"7155",
	227 => X"74B8",
	228 => X"77AD",
	229 => X"7A33",
	230 => X"7C46",
	231 => X"7DE6",
	232 => X"7F10",
	233 => X"7FC3",
	234 => X"7FFF",
	235 => X"7FC3",
	236 => X"7F10",
	237 => X"7DE6",
	238 => X"7C46",
	239 => X"7A33",
	240 => X"77AD",
	241 => X"74B8",
	242 => X"7155",
	243 => X"6D89",
	244 => X"6956",
	245 => X"64C1",
	246 => X"5FCE",
	247 => X"5A81",
	others => X"0000"
);

CONSTANT E4: hex := (
	000 => X"0000",
	001 => X"0833",
	002 => X"105E",
	003 => X"1877",
	004 => X"2077",
	005 => X"2855",
	006 => X"3008",
	007 => X"3789",
	008 => X"3ECF",
	009 => X"45D3",
	010 => X"4C8E",
	011 => X"52F8",
	012 => X"590B",
	013 => X"5EC0",
	014 => X"6412",
	015 => X"68FA",
	016 => X"6D74",
	017 => X"717B",
	018 => X"750A",
	019 => X"781E",
	020 => X"7AB4",
	021 => X"7CC9",
	022 => X"7E5A",
	023 => X"7F67",
	024 => X"7FEE",
	025 => X"7FEE",
	026 => X"7F67",
	027 => X"7E5A",
	028 => X"7CC9",
	029 => X"7AB4",
	030 => X"781E",
	031 => X"750A",
	032 => X"717B",
	033 => X"6D74",
	034 => X"68FA",
	035 => X"6412",
	036 => X"5EC0",
	037 => X"590B",
	038 => X"52F8",
	039 => X"4C8E",
	040 => X"45D3",
	041 => X"3ECF",
	042 => X"3789",
	043 => X"3008",
	044 => X"2855",
	045 => X"2077",
	046 => X"1877",
	047 => X"105E",
	048 => X"0833",
	049 => X"0000",
	050 => X"F7CB",
	051 => X"EFA0",
	052 => X"E787",
	053 => X"DF87",
	054 => X"D7A9",
	055 => X"CFF6",
	056 => X"C875",
	057 => X"C12F",
	058 => X"BA2B",
	059 => X"B370",
	060 => X"AD06",
	061 => X"A6F3",
	062 => X"A13E",
	063 => X"9BEC",
	064 => X"9704",
	065 => X"928A",
	066 => X"8E83",
	067 => X"8AF4",
	068 => X"87E0",
	069 => X"854A",
	070 => X"8335",
	071 => X"81A4",
	072 => X"8097",
	073 => X"8010",
	074 => X"8010",
	075 => X"8097",
	076 => X"81A4",
	077 => X"8335",
	078 => X"854A",
	079 => X"87E0",
	080 => X"8AF4",
	081 => X"8E83",
	082 => X"928A",
	083 => X"9704",
	084 => X"9BEC",
	085 => X"A13E",
	086 => X"A6F3",
	087 => X"AD06",
	088 => X"B370",
	089 => X"BA2B",
	090 => X"C12F",
	091 => X"C875",
	092 => X"CFF6",
	093 => X"D7A9",
	094 => X"DF87",
	095 => X"E787",
	096 => X"EFA0",
	097 => X"F7CB",
	098 => X"0000",
	099 => X"0833",
	100 => X"105E",
	101 => X"1877",
	102 => X"2077",
	103 => X"2855",
	104 => X"3008",
	105 => X"3789",
	106 => X"3ECF",
	107 => X"45D3",
	108 => X"4C8E",
	109 => X"52F8",
	110 => X"590B",
	111 => X"5EC0",
	112 => X"6412",
	113 => X"68FA",
	114 => X"6D74",
	115 => X"717B",
	116 => X"750A",
	117 => X"781E",
	118 => X"7AB4",
	119 => X"7CC9",
	120 => X"7E5A",
	121 => X"7F67",
	122 => X"7FEE",
	123 => X"7FEE",
	124 => X"7F67",
	125 => X"7E5A",
	126 => X"7CC9",
	127 => X"7AB4",
	128 => X"781E",
	129 => X"750A",
	130 => X"717B",
	131 => X"6D74",
	132 => X"68FA",
	133 => X"6412",
	134 => X"5EC0",
	135 => X"590B",
	136 => X"52F8",
	137 => X"4C8E",
	138 => X"45D3",
	139 => X"3ECF",
	140 => X"3789",
	141 => X"3008",
	142 => X"2855",
	143 => X"2077",
	144 => X"1877",
	145 => X"105E",
	146 => X"0833",
	147 => X"FFFE",
	148 => X"F7CB",
	149 => X"EFA0",
	150 => X"E787",
	151 => X"DF87",
	152 => X"D7A9",
	153 => X"CFF6",
	154 => X"C875",
	155 => X"C12F",
	156 => X"BA2B",
	157 => X"B370",
	158 => X"AD06",
	159 => X"A6F3",
	160 => X"A13E",
	161 => X"9BEC",
	162 => X"9704",
	163 => X"928A",
	164 => X"8E83",
	165 => X"8AF4",
	166 => X"87E0",
	167 => X"854A",
	168 => X"8335",
	169 => X"81A4",
	170 => X"8097",
	171 => X"8010",
	172 => X"8010",
	173 => X"8097",
	174 => X"81A4",
	175 => X"8335",
	176 => X"854A",
	177 => X"87E0",
	178 => X"8AF4",
	179 => X"8E83",
	180 => X"928A",
	181 => X"9704",
	182 => X"9BEC",
	183 => X"A13E",
	184 => X"A6F3",
	185 => X"AD06",
	186 => X"B370",
	187 => X"BA2B",
	188 => X"C12F",
	189 => X"C875",
	190 => X"CFF6",
	191 => X"D7A9",
	192 => X"DF87",
	193 => X"E787",
	194 => X"EFA0",
	195 => X"F7CB",
	196 => X"FFFE",
	197 => X"0833",
	198 => X"105E",
	199 => X"1877",
	200 => X"2077",
	201 => X"2855",
	202 => X"3008",
	203 => X"3789",
	204 => X"3ECF",
	205 => X"45D3",
	206 => X"4C8E",
	207 => X"52F8",
	208 => X"590B",
	209 => X"5EC0",
	210 => X"6412",
	211 => X"68FA",
	212 => X"6D74",
	213 => X"717B",
	214 => X"750A",
	215 => X"781E",
	216 => X"7AB4",
	217 => X"7CC9",
	218 => X"7E5A",
	219 => X"7F67",
	220 => X"7FEE",
	221 => X"7FEE",
	222 => X"7F67",
	223 => X"7E5A",
	224 => X"7CC9",
	225 => X"7AB4",
	226 => X"781E",
	227 => X"750A",
	228 => X"717B",
	229 => X"6D74",
	230 => X"68FA",
	231 => X"6412",
	232 => X"5EC0",
	233 => X"590B",
	234 => X"52F8",
	235 => X"4C8E",
	236 => X"45D3",
	237 => X"3ECF",
	238 => X"3789",
	239 => X"3008",
	240 => X"2855",
	241 => X"2077",
	242 => X"1877",
	243 => X"105E",
	244 => X"0833",
	245 => X"0000",
	246 => X"F7CB",
	247 => X"EFA0",
	others => X"0000"
);

CONSTANT F4: hex := (
	000 => X"0000",
	001 => X"08A4",
	002 => X"113E",
	003 => X"19C3",
	004 => X"222B",
	005 => X"2A6B",
	006 => X"3279",
	007 => X"3A4D",
	008 => X"41DC",
	009 => X"491E",
	010 => X"500B",
	011 => X"569B",
	012 => X"5CC5",
	013 => X"6283",
	014 => X"67CD",
	015 => X"6C9F",
	016 => X"70F2",
	017 => X"74C0",
	018 => X"7807",
	019 => X"7AC1",
	020 => X"7CEC",
	021 => X"7E85",
	022 => X"7F8A",
	023 => X"7FFA",
	024 => X"7FD4",
	025 => X"7F1A",
	026 => X"7DCB",
	027 => X"7BE8",
	028 => X"7976",
	029 => X"7675",
	030 => X"72EA",
	031 => X"6ED9",
	032 => X"6A46",
	033 => X"6537",
	034 => X"5FB2",
	035 => X"59BD",
	036 => X"535F",
	037 => X"4CA0",
	038 => X"4587",
	039 => X"3E1D",
	040 => X"366B",
	041 => X"2E79",
	042 => X"2651",
	043 => X"1DFC",
	044 => X"1584",
	045 => X"0CF2",
	046 => X"0452",
	047 => X"FBAC",
	048 => X"F30C",
	049 => X"EA7A",
	050 => X"E202",
	051 => X"D9AD",
	052 => X"D185",
	053 => X"C993",
	054 => X"C1E1",
	055 => X"BA77",
	056 => X"B35E",
	057 => X"AC9F",
	058 => X"A641",
	059 => X"A04C",
	060 => X"9AC7",
	061 => X"95B8",
	062 => X"9125",
	063 => X"8D14",
	064 => X"8989",
	065 => X"8688",
	066 => X"8416",
	067 => X"8233",
	068 => X"80E4",
	069 => X"802A",
	070 => X"8004",
	071 => X"8074",
	072 => X"8179",
	073 => X"8312",
	074 => X"853D",
	075 => X"87F7",
	076 => X"8B3E",
	077 => X"8F0C",
	078 => X"935F",
	079 => X"9831",
	080 => X"9D7B",
	081 => X"A339",
	082 => X"A963",
	083 => X"AFF3",
	084 => X"B6E0",
	085 => X"BE22",
	086 => X"C5B1",
	087 => X"CD85",
	088 => X"D593",
	089 => X"DDD3",
	090 => X"E63B",
	091 => X"EEC0",
	092 => X"F75A",
	093 => X"0000",
	094 => X"08A4",
	095 => X"113E",
	096 => X"19C3",
	097 => X"222B",
	098 => X"2A6B",
	099 => X"3279",
	100 => X"3A4D",
	101 => X"41DC",
	102 => X"491E",
	103 => X"500B",
	104 => X"569B",
	105 => X"5CC5",
	106 => X"6283",
	107 => X"67CD",
	108 => X"6C9F",
	109 => X"70F2",
	110 => X"74C0",
	111 => X"7807",
	112 => X"7AC1",
	113 => X"7CEC",
	114 => X"7E85",
	115 => X"7F8A",
	116 => X"7FFA",
	117 => X"7FD4",
	118 => X"7F1A",
	119 => X"7DCB",
	120 => X"7BE8",
	121 => X"7976",
	122 => X"7675",
	123 => X"72EA",
	124 => X"6ED9",
	125 => X"6A46",
	126 => X"6537",
	127 => X"5FB2",
	128 => X"59BD",
	129 => X"535F",
	130 => X"4CA0",
	131 => X"4587",
	132 => X"3E1D",
	133 => X"366B",
	134 => X"2E79",
	135 => X"2651",
	136 => X"1DFC",
	137 => X"1584",
	138 => X"0CF2",
	139 => X"0452",
	140 => X"FBAC",
	141 => X"F30C",
	142 => X"EA7A",
	143 => X"E202",
	144 => X"D9AD",
	145 => X"D185",
	146 => X"C993",
	147 => X"C1E1",
	148 => X"BA77",
	149 => X"B35E",
	150 => X"AC9F",
	151 => X"A641",
	152 => X"A04C",
	153 => X"9AC7",
	154 => X"95B8",
	155 => X"9125",
	156 => X"8D14",
	157 => X"8989",
	158 => X"8688",
	159 => X"8416",
	160 => X"8233",
	161 => X"80E4",
	162 => X"802A",
	163 => X"8004",
	164 => X"8074",
	165 => X"8179",
	166 => X"8312",
	167 => X"853D",
	168 => X"87F7",
	169 => X"8B3E",
	170 => X"8F0C",
	171 => X"935F",
	172 => X"9831",
	173 => X"9D7B",
	174 => X"A339",
	175 => X"A963",
	176 => X"AFF3",
	177 => X"B6E0",
	178 => X"BE22",
	179 => X"C5B1",
	180 => X"CD85",
	181 => X"D593",
	182 => X"DDD3",
	183 => X"E63B",
	184 => X"EEC0",
	185 => X"F75A",
	186 => X"0000",
	187 => X"08A4",
	188 => X"113E",
	189 => X"19C3",
	190 => X"222B",
	191 => X"2A6B",
	192 => X"3279",
	193 => X"3A4D",
	194 => X"41DC",
	195 => X"491E",
	196 => X"500B",
	197 => X"569B",
	198 => X"5CC5",
	199 => X"6283",
	200 => X"67CD",
	201 => X"6C9F",
	202 => X"70F2",
	203 => X"74C0",
	204 => X"7807",
	205 => X"7AC1",
	206 => X"7CEC",
	207 => X"7E85",
	208 => X"7F8A",
	209 => X"7FFA",
	210 => X"7FD4",
	211 => X"7F1A",
	212 => X"7DCB",
	213 => X"7BE8",
	214 => X"7976",
	215 => X"7675",
	216 => X"72EA",
	217 => X"6ED9",
	218 => X"6A46",
	219 => X"6537",
	220 => X"5FB2",
	221 => X"59BD",
	222 => X"535F",
	223 => X"4CA0",
	224 => X"4587",
	225 => X"3E1D",
	226 => X"366B",
	227 => X"2E79",
	228 => X"2651",
	229 => X"1DFC",
	230 => X"1584",
	231 => X"0CF2",
	232 => X"0452",
	233 => X"FBAC",
	234 => X"F30C",
	235 => X"EA7A",
	236 => X"E202",
	237 => X"D9AD",
	238 => X"D185",
	239 => X"C993",
	240 => X"C1E1",
	241 => X"BA77",
	242 => X"B35E",
	243 => X"AC9F",
	244 => X"A641",
	245 => X"A04C",
	246 => X"9AC7",
	247 => X"95B8",
	others => X"0000"
);

CONSTANT FS4: hex := (
	000 => X"0000",
	001 => X"0921",
	002 => X"1237",
	003 => X"1B35",
	004 => X"240F",
	005 => X"2CBA",
	006 => X"352B",
	007 => X"3D57",
	008 => X"4533",
	009 => X"4CB4",
	010 => X"53D1",
	011 => X"5A81",
	012 => X"60BB",
	013 => X"6677",
	014 => X"6BAD",
	015 => X"7056",
	016 => X"746D",
	017 => X"77ED",
	018 => X"7ACF",
	019 => X"7D12",
	020 => X"7EB1",
	021 => X"7FAB",
	022 => X"7FFF",
	023 => X"7FAB",
	024 => X"7EB1",
	025 => X"7D12",
	026 => X"7ACF",
	027 => X"77ED",
	028 => X"746D",
	029 => X"7056",
	030 => X"6BAD",
	031 => X"6677",
	032 => X"60BB",
	033 => X"5A81",
	034 => X"53D1",
	035 => X"4CB4",
	036 => X"4533",
	037 => X"3D57",
	038 => X"352B",
	039 => X"2CBA",
	040 => X"240F",
	041 => X"1B35",
	042 => X"1237",
	043 => X"0921",
	044 => X"FFFE",
	045 => X"F6DD",
	046 => X"EDC7",
	047 => X"E4C9",
	048 => X"DBEF",
	049 => X"D344",
	050 => X"CAD3",
	051 => X"C2A7",
	052 => X"BACB",
	053 => X"B34A",
	054 => X"AC2D",
	055 => X"A57D",
	056 => X"9F43",
	057 => X"9987",
	058 => X"9451",
	059 => X"8FA8",
	060 => X"8B91",
	061 => X"8811",
	062 => X"852F",
	063 => X"82EC",
	064 => X"814D",
	065 => X"8053",
	066 => X"8000",
	067 => X"8053",
	068 => X"814D",
	069 => X"82EC",
	070 => X"852F",
	071 => X"8811",
	072 => X"8B91",
	073 => X"8FA8",
	074 => X"9451",
	075 => X"9987",
	076 => X"9F43",
	077 => X"A57D",
	078 => X"AC2D",
	079 => X"B34A",
	080 => X"BACB",
	081 => X"C2A7",
	082 => X"CAD3",
	083 => X"D344",
	084 => X"DBEF",
	085 => X"E4C9",
	086 => X"EDC7",
	087 => X"F6DD",
	088 => X"FFFE",
	089 => X"0921",
	090 => X"1237",
	091 => X"1B35",
	092 => X"240F",
	093 => X"2CBA",
	094 => X"352B",
	095 => X"3D57",
	096 => X"4533",
	097 => X"4CB4",
	098 => X"53D1",
	099 => X"5A81",
	100 => X"60BB",
	101 => X"6677",
	102 => X"6BAD",
	103 => X"7056",
	104 => X"746D",
	105 => X"77ED",
	106 => X"7ACF",
	107 => X"7D12",
	108 => X"7EB1",
	109 => X"7FAB",
	110 => X"7FFF",
	111 => X"7FAB",
	112 => X"7EB1",
	113 => X"7D12",
	114 => X"7ACF",
	115 => X"77ED",
	116 => X"746D",
	117 => X"7056",
	118 => X"6BAD",
	119 => X"6677",
	120 => X"60BB",
	121 => X"5A81",
	122 => X"53D1",
	123 => X"4CB4",
	124 => X"4533",
	125 => X"3D57",
	126 => X"352B",
	127 => X"2CBA",
	128 => X"240F",
	129 => X"1B35",
	130 => X"1237",
	131 => X"0921",
	132 => X"0000",
	133 => X"F6DD",
	134 => X"EDC7",
	135 => X"E4C9",
	136 => X"DBEF",
	137 => X"D344",
	138 => X"CAD3",
	139 => X"C2A7",
	140 => X"BACB",
	141 => X"B34A",
	142 => X"AC2D",
	143 => X"A57D",
	144 => X"9F43",
	145 => X"9987",
	146 => X"9451",
	147 => X"8FA8",
	148 => X"8B91",
	149 => X"8811",
	150 => X"852F",
	151 => X"82EC",
	152 => X"814D",
	153 => X"8053",
	154 => X"8000",
	155 => X"8053",
	156 => X"814D",
	157 => X"82EC",
	158 => X"852F",
	159 => X"8811",
	160 => X"8B91",
	161 => X"8FA8",
	162 => X"9451",
	163 => X"9987",
	164 => X"9F43",
	165 => X"A57D",
	166 => X"AC2D",
	167 => X"B34A",
	168 => X"BACB",
	169 => X"C2A7",
	170 => X"CAD3",
	171 => X"D344",
	172 => X"DBEF",
	173 => X"E4C9",
	174 => X"EDC7",
	175 => X"F6DD",
	176 => X"0000",
	177 => X"0921",
	178 => X"1237",
	179 => X"1B35",
	180 => X"240F",
	181 => X"2CBA",
	182 => X"352B",
	183 => X"3D57",
	184 => X"4533",
	185 => X"4CB4",
	186 => X"53D1",
	187 => X"5A81",
	188 => X"60BB",
	189 => X"6677",
	190 => X"6BAD",
	191 => X"7056",
	192 => X"746D",
	193 => X"77ED",
	194 => X"7ACF",
	195 => X"7D12",
	196 => X"7EB1",
	197 => X"7FAB",
	198 => X"7FFF",
	199 => X"7FAB",
	200 => X"7EB1",
	201 => X"7D12",
	202 => X"7ACF",
	203 => X"77ED",
	204 => X"746D",
	205 => X"7056",
	206 => X"6BAD",
	207 => X"6677",
	208 => X"60BB",
	209 => X"5A81",
	210 => X"53D1",
	211 => X"4CB4",
	212 => X"4533",
	213 => X"3D57",
	214 => X"352B",
	215 => X"2CBA",
	216 => X"240F",
	217 => X"1B35",
	218 => X"1237",
	219 => X"0921",
	220 => X"FFFE",
	221 => X"F6DD",
	222 => X"EDC7",
	223 => X"E4C9",
	224 => X"DBEF",
	225 => X"D344",
	226 => X"CAD3",
	227 => X"C2A7",
	228 => X"BACB",
	229 => X"B34A",
	230 => X"AC2D",
	231 => X"A57D",
	232 => X"9F43",
	233 => X"9987",
	234 => X"9451",
	235 => X"8FA8",
	236 => X"8B91",
	237 => X"8811",
	238 => X"852F",
	239 => X"82EC",
	240 => X"814D",
	241 => X"8053",
	242 => X"8000",
	243 => X"8053",
	244 => X"814D",
	245 => X"82EC",
	246 => X"852F",
	247 => X"8811",
	others => X"0000"
);

CONSTANT G4: hex := (
	000 => X"0000",
	001 => X"09AE",
	002 => X"134E",
	003 => X"1CD1",
	004 => X"262B",
	005 => X"2F4C",
	006 => X"3828",
	007 => X"40B2",
	008 => X"48DD",
	009 => X"509D",
	010 => X"57E6",
	011 => X"5EAF",
	012 => X"64ED",
	013 => X"6A97",
	014 => X"6FA5",
	015 => X"740F",
	016 => X"77CF",
	017 => X"7ADF",
	018 => X"7D3B",
	019 => X"7EDF",
	020 => X"7FCA",
	021 => X"7FF9",
	022 => X"7F6C",
	023 => X"7E24",
	024 => X"7C24",
	025 => X"796D",
	026 => X"7605",
	027 => X"71EF",
	028 => X"6D32",
	029 => X"67D5",
	030 => X"61E0",
	031 => X"5B5B",
	032 => X"5451",
	033 => X"4CCB",
	034 => X"44D4",
	035 => X"3C78",
	036 => X"33C3",
	037 => X"2AC3",
	038 => X"2184",
	039 => X"1814",
	040 => X"0E80",
	041 => X"04D7",
	042 => X"FB27",
	043 => X"F17E",
	044 => X"E7EA",
	045 => X"DE7A",
	046 => X"D53B",
	047 => X"CC3B",
	048 => X"C386",
	049 => X"BB2A",
	050 => X"B333",
	051 => X"ABAD",
	052 => X"A4A3",
	053 => X"9E1E",
	054 => X"9829",
	055 => X"92CC",
	056 => X"8E0F",
	057 => X"89F9",
	058 => X"8691",
	059 => X"83DA",
	060 => X"81DA",
	061 => X"8092",
	062 => X"8005",
	063 => X"8034",
	064 => X"811F",
	065 => X"82C3",
	066 => X"851F",
	067 => X"882F",
	068 => X"8BEF",
	069 => X"9059",
	070 => X"9567",
	071 => X"9B11",
	072 => X"A14F",
	073 => X"A818",
	074 => X"AF61",
	075 => X"B721",
	076 => X"BF4C",
	077 => X"C7D6",
	078 => X"D0B2",
	079 => X"D9D3",
	080 => X"E32D",
	081 => X"ECB0",
	082 => X"F650",
	083 => X"FFFE",
	084 => X"09AE",
	085 => X"134E",
	086 => X"1CD1",
	087 => X"262B",
	088 => X"2F4C",
	089 => X"3828",
	090 => X"40B2",
	091 => X"48DD",
	092 => X"509D",
	093 => X"57E6",
	094 => X"5EAF",
	095 => X"64ED",
	096 => X"6A97",
	097 => X"6FA5",
	098 => X"740F",
	099 => X"77CF",
	100 => X"7ADF",
	101 => X"7D3B",
	102 => X"7EDF",
	103 => X"7FCA",
	104 => X"7FF9",
	105 => X"7F6C",
	106 => X"7E24",
	107 => X"7C24",
	108 => X"796D",
	109 => X"7605",
	110 => X"71EF",
	111 => X"6D32",
	112 => X"67D5",
	113 => X"61E0",
	114 => X"5B5B",
	115 => X"5451",
	116 => X"4CCB",
	117 => X"44D4",
	118 => X"3C78",
	119 => X"33C3",
	120 => X"2AC3",
	121 => X"2184",
	122 => X"1814",
	123 => X"0E80",
	124 => X"04D7",
	125 => X"FB27",
	126 => X"F17E",
	127 => X"E7EA",
	128 => X"DE7A",
	129 => X"D53B",
	130 => X"CC3B",
	131 => X"C386",
	132 => X"BB2A",
	133 => X"B333",
	134 => X"ABAD",
	135 => X"A4A3",
	136 => X"9E1E",
	137 => X"9829",
	138 => X"92CC",
	139 => X"8E0F",
	140 => X"89F9",
	141 => X"8691",
	142 => X"83DA",
	143 => X"81DA",
	144 => X"8092",
	145 => X"8005",
	146 => X"8034",
	147 => X"811F",
	148 => X"82C3",
	149 => X"851F",
	150 => X"882F",
	151 => X"8BEF",
	152 => X"9059",
	153 => X"9567",
	154 => X"9B11",
	155 => X"A14F",
	156 => X"A818",
	157 => X"AF61",
	158 => X"B721",
	159 => X"BF4C",
	160 => X"C7D6",
	161 => X"D0B2",
	162 => X"D9D3",
	163 => X"E32D",
	164 => X"ECB0",
	165 => X"F650",
	166 => X"0000",
	167 => X"09AE",
	168 => X"134E",
	169 => X"1CD1",
	170 => X"262B",
	171 => X"2F4C",
	172 => X"3828",
	173 => X"40B2",
	174 => X"48DD",
	175 => X"509D",
	176 => X"57E6",
	177 => X"5EAF",
	178 => X"64ED",
	179 => X"6A97",
	180 => X"6FA5",
	181 => X"740F",
	182 => X"77CF",
	183 => X"7ADF",
	184 => X"7D3B",
	185 => X"7EDF",
	186 => X"7FCA",
	187 => X"7FF9",
	188 => X"7F6C",
	189 => X"7E24",
	190 => X"7C24",
	191 => X"796D",
	192 => X"7605",
	193 => X"71EF",
	194 => X"6D32",
	195 => X"67D5",
	196 => X"61E0",
	197 => X"5B5B",
	198 => X"5451",
	199 => X"4CCB",
	200 => X"44D4",
	201 => X"3C78",
	202 => X"33C3",
	203 => X"2AC3",
	204 => X"2184",
	205 => X"1814",
	206 => X"0E80",
	207 => X"04D7",
	208 => X"FB27",
	209 => X"F17E",
	210 => X"E7EA",
	211 => X"DE7A",
	212 => X"D53B",
	213 => X"CC3B",
	214 => X"C386",
	215 => X"BB2A",
	216 => X"B333",
	217 => X"ABAD",
	218 => X"A4A3",
	219 => X"9E1E",
	220 => X"9829",
	221 => X"92CC",
	222 => X"8E0F",
	223 => X"89F9",
	224 => X"8691",
	225 => X"83DA",
	226 => X"81DA",
	227 => X"8092",
	228 => X"8005",
	229 => X"8034",
	230 => X"811F",
	231 => X"82C3",
	232 => X"851F",
	233 => X"882F",
	234 => X"8BEF",
	235 => X"9059",
	236 => X"9567",
	237 => X"9B11",
	238 => X"A14F",
	239 => X"A818",
	240 => X"AF61",
	241 => X"B721",
	242 => X"BF4C",
	243 => X"C7D6",
	244 => X"D0B2",
	245 => X"D9D3",
	246 => X"E32D",
	247 => X"ECB0",
	others => X"0000"
);

CONSTANT GS4: hex := (
	000 => X"0000",
	001 => X"0A4C",
	002 => X"1488",
	003 => X"1EA1",
	004 => X"2888",
	005 => X"322B",
	006 => X"3B7B",
	007 => X"4468",
	008 => X"4CE4",
	009 => X"54E0",
	010 => X"5C4F",
	011 => X"6325",
	012 => X"6956",
	013 => X"6ED9",
	014 => X"73A3",
	015 => X"77AD",
	016 => X"7AF1",
	017 => X"7D68",
	018 => X"7F10",
	019 => X"7FE4",
	020 => X"7FE4",
	021 => X"7F10",
	022 => X"7D68",
	023 => X"7AF1",
	024 => X"77AD",
	025 => X"73A3",
	026 => X"6ED9",
	027 => X"6956",
	028 => X"6325",
	029 => X"5C4F",
	030 => X"54E0",
	031 => X"4CE4",
	032 => X"4468",
	033 => X"3B7B",
	034 => X"322B",
	035 => X"2888",
	036 => X"1EA1",
	037 => X"1488",
	038 => X"0A4C",
	039 => X"0000",
	040 => X"F5B2",
	041 => X"EB76",
	042 => X"E15D",
	043 => X"D776",
	044 => X"CDD3",
	045 => X"C483",
	046 => X"BB96",
	047 => X"B31A",
	048 => X"AB1E",
	049 => X"A3AF",
	050 => X"9CD9",
	051 => X"96A8",
	052 => X"9125",
	053 => X"8C5B",
	054 => X"8851",
	055 => X"850D",
	056 => X"8296",
	057 => X"80EE",
	058 => X"801A",
	059 => X"801A",
	060 => X"80EE",
	061 => X"8296",
	062 => X"850D",
	063 => X"8851",
	064 => X"8C5B",
	065 => X"9125",
	066 => X"96A8",
	067 => X"9CD9",
	068 => X"A3AF",
	069 => X"AB1E",
	070 => X"B31A",
	071 => X"BB96",
	072 => X"C483",
	073 => X"CDD3",
	074 => X"D776",
	075 => X"E15D",
	076 => X"EB76",
	077 => X"F5B2",
	078 => X"0000",
	079 => X"0A4C",
	080 => X"1488",
	081 => X"1EA1",
	082 => X"2888",
	083 => X"322B",
	084 => X"3B7B",
	085 => X"4468",
	086 => X"4CE4",
	087 => X"54E0",
	088 => X"5C4F",
	089 => X"6325",
	090 => X"6956",
	091 => X"6ED9",
	092 => X"73A3",
	093 => X"77AD",
	094 => X"7AF1",
	095 => X"7D68",
	096 => X"7F10",
	097 => X"7FE4",
	098 => X"7FE4",
	099 => X"7F10",
	100 => X"7D68",
	101 => X"7AF1",
	102 => X"77AD",
	103 => X"73A3",
	104 => X"6ED9",
	105 => X"6956",
	106 => X"6325",
	107 => X"5C4F",
	108 => X"54E0",
	109 => X"4CE4",
	110 => X"4468",
	111 => X"3B7B",
	112 => X"322B",
	113 => X"2888",
	114 => X"1EA1",
	115 => X"1488",
	116 => X"0A4C",
	117 => X"FFFE",
	118 => X"F5B2",
	119 => X"EB76",
	120 => X"E15D",
	121 => X"D776",
	122 => X"CDD3",
	123 => X"C483",
	124 => X"BB96",
	125 => X"B31A",
	126 => X"AB1E",
	127 => X"A3AF",
	128 => X"9CD9",
	129 => X"96A8",
	130 => X"9125",
	131 => X"8C5B",
	132 => X"8851",
	133 => X"850D",
	134 => X"8296",
	135 => X"80EE",
	136 => X"801A",
	137 => X"801A",
	138 => X"80EE",
	139 => X"8296",
	140 => X"850D",
	141 => X"8851",
	142 => X"8C5B",
	143 => X"9125",
	144 => X"96A8",
	145 => X"9CD9",
	146 => X"A3AF",
	147 => X"AB1E",
	148 => X"B31A",
	149 => X"BB96",
	150 => X"C483",
	151 => X"CDD3",
	152 => X"D776",
	153 => X"E15D",
	154 => X"EB76",
	155 => X"F5B2",
	156 => X"0000",
	157 => X"0A4C",
	158 => X"1488",
	159 => X"1EA1",
	160 => X"2888",
	161 => X"322B",
	162 => X"3B7B",
	163 => X"4468",
	164 => X"4CE4",
	165 => X"54E0",
	166 => X"5C4F",
	167 => X"6325",
	168 => X"6956",
	169 => X"6ED9",
	170 => X"73A3",
	171 => X"77AD",
	172 => X"7AF1",
	173 => X"7D68",
	174 => X"7F10",
	175 => X"7FE4",
	176 => X"7FE4",
	177 => X"7F10",
	178 => X"7D68",
	179 => X"7AF1",
	180 => X"77AD",
	181 => X"73A3",
	182 => X"6ED9",
	183 => X"6956",
	184 => X"6325",
	185 => X"5C4F",
	186 => X"54E0",
	187 => X"4CE4",
	188 => X"4468",
	189 => X"3B7B",
	190 => X"322B",
	191 => X"2888",
	192 => X"1EA1",
	193 => X"1488",
	194 => X"0A4C",
	195 => X"FFFE",
	196 => X"F5B2",
	197 => X"EB76",
	198 => X"E15D",
	199 => X"D776",
	200 => X"CDD3",
	201 => X"C483",
	202 => X"BB96",
	203 => X"B31A",
	204 => X"AB1E",
	205 => X"A3AF",
	206 => X"9CD9",
	207 => X"96A8",
	208 => X"9125",
	209 => X"8C5B",
	210 => X"8851",
	211 => X"850D",
	212 => X"8296",
	213 => X"80EE",
	214 => X"801A",
	215 => X"801A",
	216 => X"80EE",
	217 => X"8296",
	218 => X"850D",
	219 => X"8851",
	220 => X"8C5B",
	221 => X"9125",
	222 => X"96A8",
	223 => X"9CD9",
	224 => X"A3AF",
	225 => X"AB1E",
	226 => X"B31A",
	227 => X"BB96",
	228 => X"C483",
	229 => X"CDD3",
	230 => X"D776",
	231 => X"E15D",
	232 => X"EB76",
	233 => X"F5B2",
	234 => X"0000",
	235 => X"0A4C",
	236 => X"1488",
	237 => X"1EA1",
	238 => X"2888",
	239 => X"322B",
	240 => X"3B7B",
	241 => X"4468",
	242 => X"4CE4",
	243 => X"54E0",
	244 => X"5C4F",
	245 => X"6325",
	246 => X"6956",
	247 => X"6ED9",
	others => X"0000"
);

CONSTANT A4: hex := (
	000 => X"0000",
	001 => X"0ADA",
	002 => X"15A1",
	003 => X"2040",
	004 => X"2AA3",
	005 => X"34B8",
	006 => X"3E6C",
	007 => X"47AC",
	008 => X"5068",
	009 => X"5890",
	010 => X"6015",
	011 => X"66E8",
	012 => X"6CFE",
	013 => X"724A",
	014 => X"76C4",
	015 => X"7A62",
	016 => X"7D1F",
	017 => X"7EF5",
	018 => X"7FE1",
	019 => X"7FE1",
	020 => X"7EF5",
	021 => X"7D1F",
	022 => X"7A62",
	023 => X"76C4",
	024 => X"724A",
	025 => X"6CFE",
	026 => X"66E8",
	027 => X"6015",
	028 => X"5890",
	029 => X"5068",
	030 => X"47AC",
	031 => X"3E6C",
	032 => X"34B8",
	033 => X"2AA3",
	034 => X"2040",
	035 => X"15A1",
	036 => X"0ADA",
	037 => X"FFFE",
	038 => X"F524",
	039 => X"EA5D",
	040 => X"DFBE",
	041 => X"D55B",
	042 => X"CB46",
	043 => X"C192",
	044 => X"B852",
	045 => X"AF96",
	046 => X"A76E",
	047 => X"9FE9",
	048 => X"9916",
	049 => X"9300",
	050 => X"8DB4",
	051 => X"893A",
	052 => X"859C",
	053 => X"82DF",
	054 => X"8109",
	055 => X"801D",
	056 => X"801D",
	057 => X"8109",
	058 => X"82DF",
	059 => X"859C",
	060 => X"893A",
	061 => X"8DB4",
	062 => X"9300",
	063 => X"9916",
	064 => X"9FE9",
	065 => X"A76E",
	066 => X"AF96",
	067 => X"B852",
	068 => X"C192",
	069 => X"CB46",
	070 => X"D55B",
	071 => X"DFBE",
	072 => X"EA5D",
	073 => X"F524",
	074 => X"FFFE",
	075 => X"0ADA",
	076 => X"15A1",
	077 => X"2040",
	078 => X"2AA3",
	079 => X"34B8",
	080 => X"3E6C",
	081 => X"47AC",
	082 => X"5068",
	083 => X"5890",
	084 => X"6015",
	085 => X"66E8",
	086 => X"6CFE",
	087 => X"724A",
	088 => X"76C4",
	089 => X"7A62",
	090 => X"7D1F",
	091 => X"7EF5",
	092 => X"7FE1",
	093 => X"7FE1",
	094 => X"7EF5",
	095 => X"7D1F",
	096 => X"7A62",
	097 => X"76C4",
	098 => X"724A",
	099 => X"6CFE",
	100 => X"66E8",
	101 => X"6015",
	102 => X"5890",
	103 => X"5068",
	104 => X"47AC",
	105 => X"3E6C",
	106 => X"34B8",
	107 => X"2AA3",
	108 => X"2040",
	109 => X"15A1",
	110 => X"0ADA",
	111 => X"0000",
	112 => X"F524",
	113 => X"EA5D",
	114 => X"DFBE",
	115 => X"D55B",
	116 => X"CB46",
	117 => X"C192",
	118 => X"B852",
	119 => X"AF96",
	120 => X"A76E",
	121 => X"9FE9",
	122 => X"9916",
	123 => X"9300",
	124 => X"8DB4",
	125 => X"893A",
	126 => X"859C",
	127 => X"82DF",
	128 => X"8109",
	129 => X"801D",
	130 => X"801D",
	131 => X"8109",
	132 => X"82DF",
	133 => X"859C",
	134 => X"893A",
	135 => X"8DB4",
	136 => X"9300",
	137 => X"9916",
	138 => X"9FE9",
	139 => X"A76E",
	140 => X"AF96",
	141 => X"B852",
	142 => X"C192",
	143 => X"CB46",
	144 => X"D55B",
	145 => X"DFBE",
	146 => X"EA5D",
	147 => X"F524",
	148 => X"0000",
	149 => X"0ADA",
	150 => X"15A1",
	151 => X"2040",
	152 => X"2AA3",
	153 => X"34B8",
	154 => X"3E6C",
	155 => X"47AC",
	156 => X"5068",
	157 => X"5890",
	158 => X"6015",
	159 => X"66E8",
	160 => X"6CFE",
	161 => X"724A",
	162 => X"76C4",
	163 => X"7A62",
	164 => X"7D1F",
	165 => X"7EF5",
	166 => X"7FE1",
	167 => X"7FE1",
	168 => X"7EF5",
	169 => X"7D1F",
	170 => X"7A62",
	171 => X"76C4",
	172 => X"724A",
	173 => X"6CFE",
	174 => X"66E8",
	175 => X"6015",
	176 => X"5890",
	177 => X"5068",
	178 => X"47AC",
	179 => X"3E6C",
	180 => X"34B8",
	181 => X"2AA3",
	182 => X"2040",
	183 => X"15A1",
	184 => X"0ADA",
	185 => X"FFFE",
	186 => X"F524",
	187 => X"EA5D",
	188 => X"DFBE",
	189 => X"D55B",
	190 => X"CB46",
	191 => X"C192",
	192 => X"B852",
	193 => X"AF96",
	194 => X"A76E",
	195 => X"9FE9",
	196 => X"9916",
	197 => X"9300",
	198 => X"8DB4",
	199 => X"893A",
	200 => X"859C",
	201 => X"82DF",
	202 => X"8109",
	203 => X"801D",
	204 => X"801D",
	205 => X"8109",
	206 => X"82DF",
	207 => X"859C",
	208 => X"893A",
	209 => X"8DB4",
	210 => X"9300",
	211 => X"9916",
	212 => X"9FE9",
	213 => X"A76E",
	214 => X"AF96",
	215 => X"B852",
	216 => X"C192",
	217 => X"CB46",
	218 => X"D55B",
	219 => X"DFBE",
	220 => X"EA5D",
	221 => X"F524",
	222 => X"0000",
	223 => X"0ADA",
	224 => X"15A1",
	225 => X"2040",
	226 => X"2AA3",
	227 => X"34B8",
	228 => X"3E6C",
	229 => X"47AC",
	230 => X"5068",
	231 => X"5890",
	232 => X"6015",
	233 => X"66E8",
	234 => X"6CFE",
	235 => X"724A",
	236 => X"76C4",
	237 => X"7A62",
	238 => X"7D1F",
	239 => X"7EF5",
	240 => X"7FE1",
	241 => X"7FE1",
	242 => X"7EF5",
	243 => X"7D1F",
	244 => X"7A62",
	245 => X"76C4",
	246 => X"724A",
	247 => X"6CFE",
	others => X"0000"
);

CONSTANT AS4: hex := (
	000 => X"0000",
	001 => X"0B79",
	002 => X"16DA",
	003 => X"220D",
	004 => X"2CF9",
	005 => X"3789",
	006 => X"41A6",
	007 => X"4B3B",
	008 => X"5436",
	009 => X"5C83",
	010 => X"6412",
	011 => X"6AD2",
	012 => X"70B6",
	013 => X"75B2",
	014 => X"79BB",
	015 => X"7CC9",
	016 => X"7ED6",
	017 => X"7FDE",
	018 => X"7FDE",
	019 => X"7ED6",
	020 => X"7CC9",
	021 => X"79BB",
	022 => X"75B2",
	023 => X"70B6",
	024 => X"6AD2",
	025 => X"6412",
	026 => X"5C83",
	027 => X"5436",
	028 => X"4B3B",
	029 => X"41A6",
	030 => X"3789",
	031 => X"2CF9",
	032 => X"220D",
	033 => X"16DA",
	034 => X"0B79",
	035 => X"0000",
	036 => X"F485",
	037 => X"E924",
	038 => X"DDF1",
	039 => X"D305",
	040 => X"C875",
	041 => X"BE58",
	042 => X"B4C3",
	043 => X"ABC8",
	044 => X"A37B",
	045 => X"9BEC",
	046 => X"952C",
	047 => X"8F48",
	048 => X"8A4C",
	049 => X"8643",
	050 => X"8335",
	051 => X"8128",
	052 => X"8020",
	053 => X"8020",
	054 => X"8128",
	055 => X"8335",
	056 => X"8643",
	057 => X"8A4C",
	058 => X"8F48",
	059 => X"952C",
	060 => X"9BEC",
	061 => X"A37B",
	062 => X"ABC8",
	063 => X"B4C3",
	064 => X"BE58",
	065 => X"C875",
	066 => X"D305",
	067 => X"DDF1",
	068 => X"E924",
	069 => X"F485",
	070 => X"0000",
	071 => X"0B79",
	072 => X"16DA",
	073 => X"220D",
	074 => X"2CF9",
	075 => X"3789",
	076 => X"41A6",
	077 => X"4B3B",
	078 => X"5436",
	079 => X"5C83",
	080 => X"6412",
	081 => X"6AD2",
	082 => X"70B6",
	083 => X"75B2",
	084 => X"79BB",
	085 => X"7CC9",
	086 => X"7ED6",
	087 => X"7FDE",
	088 => X"7FDE",
	089 => X"7ED6",
	090 => X"7CC9",
	091 => X"79BB",
	092 => X"75B2",
	093 => X"70B6",
	094 => X"6AD2",
	095 => X"6412",
	096 => X"5C83",
	097 => X"5436",
	098 => X"4B3B",
	099 => X"41A6",
	100 => X"3789",
	101 => X"2CF9",
	102 => X"220D",
	103 => X"16DA",
	104 => X"0B79",
	105 => X"FFFE",
	106 => X"F485",
	107 => X"E924",
	108 => X"DDF1",
	109 => X"D305",
	110 => X"C875",
	111 => X"BE58",
	112 => X"B4C3",
	113 => X"ABC8",
	114 => X"A37B",
	115 => X"9BEC",
	116 => X"952C",
	117 => X"8F48",
	118 => X"8A4C",
	119 => X"8643",
	120 => X"8335",
	121 => X"8128",
	122 => X"8020",
	123 => X"8020",
	124 => X"8128",
	125 => X"8335",
	126 => X"8643",
	127 => X"8A4C",
	128 => X"8F48",
	129 => X"952C",
	130 => X"9BEC",
	131 => X"A37B",
	132 => X"ABC8",
	133 => X"B4C3",
	134 => X"BE58",
	135 => X"C875",
	136 => X"D305",
	137 => X"DDF1",
	138 => X"E924",
	139 => X"F485",
	140 => X"FFFE",
	141 => X"0B79",
	142 => X"16DA",
	143 => X"220D",
	144 => X"2CF9",
	145 => X"3789",
	146 => X"41A6",
	147 => X"4B3B",
	148 => X"5436",
	149 => X"5C83",
	150 => X"6412",
	151 => X"6AD2",
	152 => X"70B6",
	153 => X"75B2",
	154 => X"79BB",
	155 => X"7CC9",
	156 => X"7ED6",
	157 => X"7FDE",
	158 => X"7FDE",
	159 => X"7ED6",
	160 => X"7CC9",
	161 => X"79BB",
	162 => X"75B2",
	163 => X"70B6",
	164 => X"6AD2",
	165 => X"6412",
	166 => X"5C83",
	167 => X"5436",
	168 => X"4B3B",
	169 => X"41A6",
	170 => X"3789",
	171 => X"2CF9",
	172 => X"220D",
	173 => X"16DA",
	174 => X"0B79",
	175 => X"0000",
	176 => X"F485",
	177 => X"E924",
	178 => X"DDF1",
	179 => X"D305",
	180 => X"C875",
	181 => X"BE58",
	182 => X"B4C3",
	183 => X"ABC8",
	184 => X"A37B",
	185 => X"9BEC",
	186 => X"952C",
	187 => X"8F48",
	188 => X"8A4C",
	189 => X"8643",
	190 => X"8335",
	191 => X"8128",
	192 => X"8020",
	193 => X"8020",
	194 => X"8128",
	195 => X"8335",
	196 => X"8643",
	197 => X"8A4C",
	198 => X"8F48",
	199 => X"952C",
	200 => X"9BEC",
	201 => X"A37B",
	202 => X"ABC8",
	203 => X"B4C3",
	204 => X"BE58",
	205 => X"C875",
	206 => X"D305",
	207 => X"DDF1",
	208 => X"E924",
	209 => X"F485",
	210 => X"FFFE",
	211 => X"0B79",
	212 => X"16DA",
	213 => X"220D",
	214 => X"2CF9",
	215 => X"3789",
	216 => X"41A6",
	217 => X"4B3B",
	218 => X"5436",
	219 => X"5C83",
	220 => X"6412",
	221 => X"6AD2",
	222 => X"70B6",
	223 => X"75B2",
	224 => X"79BB",
	225 => X"7CC9",
	226 => X"7ED6",
	227 => X"7FDE",
	228 => X"7FDE",
	229 => X"7ED6",
	230 => X"7CC9",
	231 => X"79BB",
	232 => X"75B2",
	233 => X"70B6",
	234 => X"6AD2",
	235 => X"6412",
	236 => X"5C83",
	237 => X"5436",
	238 => X"4B3B",
	239 => X"41A6",
	240 => X"3789",
	241 => X"2CF9",
	242 => X"220D",
	243 => X"16DA",
	244 => X"0B79",
	245 => X"0000",
	246 => X"F485",
	247 => X"E924",
	others => X"0000"
);

CONSTANT B4: hex := (
	000 => X"0000",
	001 => X"0C2A",
	002 => X"1839",
	003 => X"240F",
	004 => X"2F92",
	005 => X"3AA6",
	006 => X"4533",
	007 => X"4F1F",
	008 => X"5853",
	009 => X"60BB",
	010 => X"6843",
	011 => X"6ED9",
	012 => X"746D",
	013 => X"78F4",
	014 => X"7C63",
	015 => X"7EB1",
	016 => X"7FD9",
	017 => X"7FD9",
	018 => X"7EB1",
	019 => X"7C63",
	020 => X"78F4",
	021 => X"746D",
	022 => X"6ED9",
	023 => X"6843",
	024 => X"60BB",
	025 => X"5853",
	026 => X"4F1F",
	027 => X"4533",
	028 => X"3AA6",
	029 => X"2F92",
	030 => X"240F",
	031 => X"1839",
	032 => X"0C2A",
	033 => X"FFFE",
	034 => X"F3D4",
	035 => X"E7C5",
	036 => X"DBEF",
	037 => X"D06C",
	038 => X"C558",
	039 => X"BACB",
	040 => X"B0DF",
	041 => X"A7AB",
	042 => X"9F43",
	043 => X"97BB",
	044 => X"9125",
	045 => X"8B91",
	046 => X"870A",
	047 => X"839B",
	048 => X"814D",
	049 => X"8025",
	050 => X"8025",
	051 => X"814D",
	052 => X"839B",
	053 => X"870A",
	054 => X"8B91",
	055 => X"9125",
	056 => X"97BB",
	057 => X"9F43",
	058 => X"A7AB",
	059 => X"B0DF",
	060 => X"BACB",
	061 => X"C558",
	062 => X"D06C",
	063 => X"DBEF",
	064 => X"E7C5",
	065 => X"F3D4",
	066 => X"FFFE",
	067 => X"0C2A",
	068 => X"1839",
	069 => X"240F",
	070 => X"2F92",
	071 => X"3AA6",
	072 => X"4533",
	073 => X"4F1F",
	074 => X"5853",
	075 => X"60BB",
	076 => X"6843",
	077 => X"6ED9",
	078 => X"746D",
	079 => X"78F4",
	080 => X"7C63",
	081 => X"7EB1",
	082 => X"7FD9",
	083 => X"7FD9",
	084 => X"7EB1",
	085 => X"7C63",
	086 => X"78F4",
	087 => X"746D",
	088 => X"6ED9",
	089 => X"6843",
	090 => X"60BB",
	091 => X"5853",
	092 => X"4F1F",
	093 => X"4533",
	094 => X"3AA6",
	095 => X"2F92",
	096 => X"240F",
	097 => X"1839",
	098 => X"0C2A",
	099 => X"0000",
	100 => X"F3D4",
	101 => X"E7C5",
	102 => X"DBEF",
	103 => X"D06C",
	104 => X"C558",
	105 => X"BACB",
	106 => X"B0DF",
	107 => X"A7AB",
	108 => X"9F43",
	109 => X"97BB",
	110 => X"9125",
	111 => X"8B91",
	112 => X"870A",
	113 => X"839B",
	114 => X"814D",
	115 => X"8025",
	116 => X"8025",
	117 => X"814D",
	118 => X"839B",
	119 => X"870A",
	120 => X"8B91",
	121 => X"9125",
	122 => X"97BB",
	123 => X"9F43",
	124 => X"A7AB",
	125 => X"B0DF",
	126 => X"BACB",
	127 => X"C558",
	128 => X"D06C",
	129 => X"DBEF",
	130 => X"E7C5",
	131 => X"F3D4",
	132 => X"0000",
	133 => X"0C2A",
	134 => X"1839",
	135 => X"240F",
	136 => X"2F92",
	137 => X"3AA6",
	138 => X"4533",
	139 => X"4F1F",
	140 => X"5853",
	141 => X"60BB",
	142 => X"6843",
	143 => X"6ED9",
	144 => X"746D",
	145 => X"78F4",
	146 => X"7C63",
	147 => X"7EB1",
	148 => X"7FD9",
	149 => X"7FD9",
	150 => X"7EB1",
	151 => X"7C63",
	152 => X"78F4",
	153 => X"746D",
	154 => X"6ED9",
	155 => X"6843",
	156 => X"60BB",
	157 => X"5853",
	158 => X"4F1F",
	159 => X"4533",
	160 => X"3AA6",
	161 => X"2F92",
	162 => X"240F",
	163 => X"1839",
	164 => X"0C2A",
	165 => X"FFFE",
	166 => X"F3D4",
	167 => X"E7C5",
	168 => X"DBEF",
	169 => X"D06C",
	170 => X"C558",
	171 => X"BACB",
	172 => X"B0DF",
	173 => X"A7AB",
	174 => X"9F43",
	175 => X"97BB",
	176 => X"9125",
	177 => X"8B91",
	178 => X"870A",
	179 => X"839B",
	180 => X"814D",
	181 => X"8025",
	182 => X"8025",
	183 => X"814D",
	184 => X"839B",
	185 => X"870A",
	186 => X"8B91",
	187 => X"9125",
	188 => X"97BB",
	189 => X"9F43",
	190 => X"A7AB",
	191 => X"B0DF",
	192 => X"BACB",
	193 => X"C558",
	194 => X"D06C",
	195 => X"DBEF",
	196 => X"E7C5",
	197 => X"F3D4",
	198 => X"0000",
	199 => X"0C2A",
	200 => X"1839",
	201 => X"240F",
	202 => X"2F92",
	203 => X"3AA6",
	204 => X"4533",
	205 => X"4F1F",
	206 => X"5853",
	207 => X"60BB",
	208 => X"6843",
	209 => X"6ED9",
	210 => X"746D",
	211 => X"78F4",
	212 => X"7C63",
	213 => X"7EB1",
	214 => X"7FD9",
	215 => X"7FD9",
	216 => X"7EB1",
	217 => X"7C63",
	218 => X"78F4",
	219 => X"746D",
	220 => X"6ED9",
	221 => X"6843",
	222 => X"60BB",
	223 => X"5853",
	224 => X"4F1F",
	225 => X"4533",
	226 => X"3AA6",
	227 => X"2F92",
	228 => X"240F",
	229 => X"1839",
	230 => X"0C2A",
	231 => X"FFFE",
	232 => X"F3D4",
	233 => X"E7C5",
	234 => X"DBEF",
	235 => X"D06C",
	236 => X"C558",
	237 => X"BACB",
	238 => X"B0DF",
	239 => X"A7AB",
	240 => X"9F43",
	241 => X"97BB",
	242 => X"9125",
	243 => X"8B91",
	244 => X"870A",
	245 => X"839B",
	246 => X"814D",
	247 => X"8025",
	others => X"0000"
);

CONSTANT C5: hex := (
	000 => X"0000",
	001 => X"0CF2",
	002 => X"19C3",
	003 => X"2651",
	004 => X"3279",
	005 => X"3E1D",
	006 => X"491E",
	007 => X"535F",
	008 => X"5CC5",
	009 => X"6537",
	010 => X"6C9F",
	011 => X"72EA",
	012 => X"7807",
	013 => X"7BE8",
	014 => X"7E85",
	015 => X"7FD4",
	016 => X"7FD4",
	017 => X"7E85",
	018 => X"7BE8",
	019 => X"7807",
	020 => X"72EA",
	021 => X"6C9F",
	022 => X"6537",
	023 => X"5CC5",
	024 => X"535F",
	025 => X"491E",
	026 => X"3E1D",
	027 => X"3279",
	028 => X"2651",
	029 => X"19C3",
	030 => X"0CF2",
	031 => X"FFFE",
	032 => X"F30C",
	033 => X"E63B",
	034 => X"D9AD",
	035 => X"CD85",
	036 => X"C1E1",
	037 => X"B6E0",
	038 => X"AC9F",
	039 => X"A339",
	040 => X"9AC7",
	041 => X"935F",
	042 => X"8D14",
	043 => X"87F7",
	044 => X"8416",
	045 => X"8179",
	046 => X"802A",
	047 => X"802A",
	048 => X"8179",
	049 => X"8416",
	050 => X"87F7",
	051 => X"8D14",
	052 => X"935F",
	053 => X"9AC7",
	054 => X"A339",
	055 => X"AC9F",
	056 => X"B6E0",
	057 => X"C1E1",
	058 => X"CD85",
	059 => X"D9AD",
	060 => X"E63B",
	061 => X"F30C",
	062 => X"0000",
	063 => X"0CF2",
	064 => X"19C3",
	065 => X"2651",
	066 => X"3279",
	067 => X"3E1D",
	068 => X"491E",
	069 => X"535F",
	070 => X"5CC5",
	071 => X"6537",
	072 => X"6C9F",
	073 => X"72EA",
	074 => X"7807",
	075 => X"7BE8",
	076 => X"7E85",
	077 => X"7FD4",
	078 => X"7FD4",
	079 => X"7E85",
	080 => X"7BE8",
	081 => X"7807",
	082 => X"72EA",
	083 => X"6C9F",
	084 => X"6537",
	085 => X"5CC5",
	086 => X"535F",
	087 => X"491E",
	088 => X"3E1D",
	089 => X"3279",
	090 => X"2651",
	091 => X"19C3",
	092 => X"0CF2",
	093 => X"FFFE",
	094 => X"F30C",
	095 => X"E63B",
	096 => X"D9AD",
	097 => X"CD85",
	098 => X"C1E1",
	099 => X"B6E0",
	100 => X"AC9F",
	101 => X"A339",
	102 => X"9AC7",
	103 => X"935F",
	104 => X"8D14",
	105 => X"87F7",
	106 => X"8416",
	107 => X"8179",
	108 => X"802A",
	109 => X"802A",
	110 => X"8179",
	111 => X"8416",
	112 => X"87F7",
	113 => X"8D14",
	114 => X"935F",
	115 => X"9AC7",
	116 => X"A339",
	117 => X"AC9F",
	118 => X"B6E0",
	119 => X"C1E1",
	120 => X"CD85",
	121 => X"D9AD",
	122 => X"E63B",
	123 => X"F30C",
	124 => X"FFFE",
	125 => X"0CF2",
	126 => X"19C3",
	127 => X"2651",
	128 => X"3279",
	129 => X"3E1D",
	130 => X"491E",
	131 => X"535F",
	132 => X"5CC5",
	133 => X"6537",
	134 => X"6C9F",
	135 => X"72EA",
	136 => X"7807",
	137 => X"7BE8",
	138 => X"7E85",
	139 => X"7FD4",
	140 => X"7FD4",
	141 => X"7E85",
	142 => X"7BE8",
	143 => X"7807",
	144 => X"72EA",
	145 => X"6C9F",
	146 => X"6537",
	147 => X"5CC5",
	148 => X"535F",
	149 => X"491E",
	150 => X"3E1D",
	151 => X"3279",
	152 => X"2651",
	153 => X"19C3",
	154 => X"0CF2",
	155 => X"0000",
	156 => X"F30C",
	157 => X"E63B",
	158 => X"D9AD",
	159 => X"CD85",
	160 => X"C1E1",
	161 => X"B6E0",
	162 => X"AC9F",
	163 => X"A339",
	164 => X"9AC7",
	165 => X"935F",
	166 => X"8D14",
	167 => X"87F7",
	168 => X"8416",
	169 => X"8179",
	170 => X"802A",
	171 => X"802A",
	172 => X"8179",
	173 => X"8416",
	174 => X"87F7",
	175 => X"8D14",
	176 => X"935F",
	177 => X"9AC7",
	178 => X"A339",
	179 => X"AC9F",
	180 => X"B6E0",
	181 => X"C1E1",
	182 => X"CD85",
	183 => X"D9AD",
	184 => X"E63B",
	185 => X"F30C",
	186 => X"FFFE",
	187 => X"0CF2",
	188 => X"19C3",
	189 => X"2651",
	190 => X"3279",
	191 => X"3E1D",
	192 => X"491E",
	193 => X"535F",
	194 => X"5CC5",
	195 => X"6537",
	196 => X"6C9F",
	197 => X"72EA",
	198 => X"7807",
	199 => X"7BE8",
	200 => X"7E85",
	201 => X"7FD4",
	202 => X"7FD4",
	203 => X"7E85",
	204 => X"7BE8",
	205 => X"7807",
	206 => X"72EA",
	207 => X"6C9F",
	208 => X"6537",
	209 => X"5CC5",
	210 => X"535F",
	211 => X"491E",
	212 => X"3E1D",
	213 => X"3279",
	214 => X"2651",
	215 => X"19C3",
	216 => X"0CF2",
	217 => X"0000",
	218 => X"F30C",
	219 => X"E63B",
	220 => X"D9AD",
	221 => X"CD85",
	222 => X"C1E1",
	223 => X"B6E0",
	224 => X"AC9F",
	225 => X"A339",
	226 => X"9AC7",
	227 => X"935F",
	228 => X"8D14",
	229 => X"87F7",
	230 => X"8416",
	231 => X"8179",
	232 => X"802A",
	233 => X"802A",
	234 => X"8179",
	235 => X"8416",
	236 => X"87F7",
	237 => X"8D14",
	238 => X"935F",
	239 => X"9AC7",
	240 => X"A339",
	241 => X"AC9F",
	242 => X"B6E0",
	243 => X"C1E1",
	244 => X"CD85",
	245 => X"D9AD",
	246 => X"E63B",
	247 => X"F30C",
	others => X"0000"
);

CONSTANT CS5: hex := (
	000 => X"0000",
	001 => X"0D9A",
	002 => X"1B0E",
	003 => X"2833",
	004 => X"34E3",
	005 => X"40FA",
	006 => X"4C55",
	007 => X"56D2",
	008 => X"6053",
	009 => X"68BD",
	010 => X"6FF7",
	011 => X"75EC",
	012 => X"7A8B",
	013 => X"7DC7",
	014 => X"7F96",
	015 => X"7FF3",
	016 => X"7EDD",
	017 => X"7C56",
	018 => X"7867",
	019 => X"731B",
	020 => X"6C81",
	021 => X"64AC",
	022 => X"5BB4",
	023 => X"51B1",
	024 => X"46C1",
	025 => X"3B04",
	026 => X"2E9C",
	027 => X"21AD",
	028 => X"145C",
	029 => X"06CF",
	030 => X"F92F",
	031 => X"EBA2",
	032 => X"DE51",
	033 => X"D162",
	034 => X"C4FA",
	035 => X"B93D",
	036 => X"AE4D",
	037 => X"A44A",
	038 => X"9B52",
	039 => X"937D",
	040 => X"8CE3",
	041 => X"8797",
	042 => X"83A8",
	043 => X"8121",
	044 => X"800B",
	045 => X"8068",
	046 => X"8237",
	047 => X"8573",
	048 => X"8A12",
	049 => X"9007",
	050 => X"9741",
	051 => X"9FAB",
	052 => X"A92C",
	053 => X"B3A9",
	054 => X"BF04",
	055 => X"CB1B",
	056 => X"D7CB",
	057 => X"E4F0",
	058 => X"F264",
	059 => X"0000",
	060 => X"0D9A",
	061 => X"1B0E",
	062 => X"2833",
	063 => X"34E3",
	064 => X"40FA",
	065 => X"4C55",
	066 => X"56D2",
	067 => X"6053",
	068 => X"68BD",
	069 => X"6FF7",
	070 => X"75EC",
	071 => X"7A8B",
	072 => X"7DC7",
	073 => X"7F96",
	074 => X"7FF3",
	075 => X"7EDD",
	076 => X"7C56",
	077 => X"7867",
	078 => X"731B",
	079 => X"6C81",
	080 => X"64AC",
	081 => X"5BB4",
	082 => X"51B1",
	083 => X"46C1",
	084 => X"3B04",
	085 => X"2E9C",
	086 => X"21AD",
	087 => X"145C",
	088 => X"06CF",
	089 => X"F92F",
	090 => X"EBA2",
	091 => X"DE51",
	092 => X"D162",
	093 => X"C4FA",
	094 => X"B93D",
	095 => X"AE4D",
	096 => X"A44A",
	097 => X"9B52",
	098 => X"937D",
	099 => X"8CE3",
	100 => X"8797",
	101 => X"83A8",
	102 => X"8121",
	103 => X"800B",
	104 => X"8068",
	105 => X"8237",
	106 => X"8573",
	107 => X"8A12",
	108 => X"9007",
	109 => X"9741",
	110 => X"9FAB",
	111 => X"A92C",
	112 => X"B3A9",
	113 => X"BF04",
	114 => X"CB1B",
	115 => X"D7CB",
	116 => X"E4F0",
	117 => X"F264",
	118 => X"0000",
	119 => X"0D9A",
	120 => X"1B0E",
	121 => X"2833",
	122 => X"34E3",
	123 => X"40FA",
	124 => X"4C55",
	125 => X"56D2",
	126 => X"6053",
	127 => X"68BD",
	128 => X"6FF7",
	129 => X"75EC",
	130 => X"7A8B",
	131 => X"7DC7",
	132 => X"7F96",
	133 => X"7FF3",
	134 => X"7EDD",
	135 => X"7C56",
	136 => X"7867",
	137 => X"731B",
	138 => X"6C81",
	139 => X"64AC",
	140 => X"5BB4",
	141 => X"51B1",
	142 => X"46C1",
	143 => X"3B04",
	144 => X"2E9C",
	145 => X"21AD",
	146 => X"145C",
	147 => X"06CF",
	148 => X"F92F",
	149 => X"EBA2",
	150 => X"DE51",
	151 => X"D162",
	152 => X"C4FA",
	153 => X"B93D",
	154 => X"AE4D",
	155 => X"A44A",
	156 => X"9B52",
	157 => X"937D",
	158 => X"8CE3",
	159 => X"8797",
	160 => X"83A8",
	161 => X"8121",
	162 => X"800B",
	163 => X"8068",
	164 => X"8237",
	165 => X"8573",
	166 => X"8A12",
	167 => X"9007",
	168 => X"9741",
	169 => X"9FAB",
	170 => X"A92C",
	171 => X"B3A9",
	172 => X"BF04",
	173 => X"CB1B",
	174 => X"D7CB",
	175 => X"E4F0",
	176 => X"F264",
	177 => X"0000",
	178 => X"0D9A",
	179 => X"1B0E",
	180 => X"2833",
	181 => X"34E3",
	182 => X"40FA",
	183 => X"4C55",
	184 => X"56D2",
	185 => X"6053",
	186 => X"68BD",
	187 => X"6FF7",
	188 => X"75EC",
	189 => X"7A8B",
	190 => X"7DC7",
	191 => X"7F96",
	192 => X"7FF3",
	193 => X"7EDD",
	194 => X"7C56",
	195 => X"7867",
	196 => X"731B",
	197 => X"6C81",
	198 => X"64AC",
	199 => X"5BB4",
	200 => X"51B1",
	201 => X"46C1",
	202 => X"3B04",
	203 => X"2E9C",
	204 => X"21AD",
	205 => X"145C",
	206 => X"06CF",
	207 => X"F92F",
	208 => X"EBA2",
	209 => X"DE51",
	210 => X"D162",
	211 => X"C4FA",
	212 => X"B93D",
	213 => X"AE4D",
	214 => X"A44A",
	215 => X"9B52",
	216 => X"937D",
	217 => X"8CE3",
	218 => X"8797",
	219 => X"83A8",
	220 => X"8121",
	221 => X"800B",
	222 => X"8068",
	223 => X"8237",
	224 => X"8573",
	225 => X"8A12",
	226 => X"9007",
	227 => X"9741",
	228 => X"9FAB",
	229 => X"A92C",
	230 => X"B3A9",
	231 => X"BF04",
	232 => X"CB1B",
	233 => X"D7CB",
	234 => X"E4F0",
	235 => X"F264",
	236 => X"0000",
	237 => X"0D9A",
	238 => X"1B0E",
	239 => X"2833",
	240 => X"34E3",
	241 => X"40FA",
	242 => X"4C55",
	243 => X"56D2",
	244 => X"6053",
	245 => X"68BD",
	246 => X"6FF7",
	247 => X"75EC",
	others => X"0000"
);

CONSTANT D5: hex := (
	000 => X"0000",
	001 => X"0E97",
	002 => X"1CFD",
	003 => X"2B03",
	004 => X"3879",
	005 => X"4533",
	006 => X"5105",
	007 => X"5BCA",
	008 => X"655C",
	009 => X"6D9B",
	010 => X"746D",
	011 => X"79BB",
	012 => X"7D72",
	013 => X"7F86",
	014 => X"7FF1",
	015 => X"7EB1",
	016 => X"7BCA",
	017 => X"7746",
	018 => X"7134",
	019 => X"69A8",
	020 => X"60BB",
	021 => X"568C",
	022 => X"4B3B",
	023 => X"3EF0",
	024 => X"31D3",
	025 => X"240F",
	026 => X"15D3",
	027 => X"074E",
	028 => X"F8B0",
	029 => X"EA2B",
	030 => X"DBEF",
	031 => X"CE2B",
	032 => X"C10E",
	033 => X"B4C3",
	034 => X"A972",
	035 => X"9F43",
	036 => X"9656",
	037 => X"8ECA",
	038 => X"88B8",
	039 => X"8434",
	040 => X"814D",
	041 => X"800D",
	042 => X"8078",
	043 => X"828C",
	044 => X"8643",
	045 => X"8B91",
	046 => X"9263",
	047 => X"9AA2",
	048 => X"A434",
	049 => X"AEF9",
	050 => X"BACB",
	051 => X"C785",
	052 => X"D4FB",
	053 => X"E301",
	054 => X"F167",
	055 => X"FFFE",
	056 => X"0E97",
	057 => X"1CFD",
	058 => X"2B03",
	059 => X"3879",
	060 => X"4533",
	061 => X"5105",
	062 => X"5BCA",
	063 => X"655C",
	064 => X"6D9B",
	065 => X"746D",
	066 => X"79BB",
	067 => X"7D72",
	068 => X"7F86",
	069 => X"7FF1",
	070 => X"7EB1",
	071 => X"7BCA",
	072 => X"7746",
	073 => X"7134",
	074 => X"69A8",
	075 => X"60BB",
	076 => X"568C",
	077 => X"4B3B",
	078 => X"3EF0",
	079 => X"31D3",
	080 => X"240F",
	081 => X"15D3",
	082 => X"074E",
	083 => X"F8B0",
	084 => X"EA2B",
	085 => X"DBEF",
	086 => X"CE2B",
	087 => X"C10E",
	088 => X"B4C3",
	089 => X"A972",
	090 => X"9F43",
	091 => X"9656",
	092 => X"8ECA",
	093 => X"88B8",
	094 => X"8434",
	095 => X"814D",
	096 => X"800D",
	097 => X"8078",
	098 => X"828C",
	099 => X"8643",
	100 => X"8B91",
	101 => X"9263",
	102 => X"9AA2",
	103 => X"A434",
	104 => X"AEF9",
	105 => X"BACB",
	106 => X"C785",
	107 => X"D4FB",
	108 => X"E301",
	109 => X"F167",
	110 => X"FFFE",
	111 => X"0E97",
	112 => X"1CFD",
	113 => X"2B03",
	114 => X"3879",
	115 => X"4533",
	116 => X"5105",
	117 => X"5BCA",
	118 => X"655C",
	119 => X"6D9B",
	120 => X"746D",
	121 => X"79BB",
	122 => X"7D72",
	123 => X"7F86",
	124 => X"7FF1",
	125 => X"7EB1",
	126 => X"7BCA",
	127 => X"7746",
	128 => X"7134",
	129 => X"69A8",
	130 => X"60BB",
	131 => X"568C",
	132 => X"4B3B",
	133 => X"3EF0",
	134 => X"31D3",
	135 => X"240F",
	136 => X"15D3",
	137 => X"074E",
	138 => X"F8B0",
	139 => X"EA2B",
	140 => X"DBEF",
	141 => X"CE2B",
	142 => X"C10E",
	143 => X"B4C3",
	144 => X"A972",
	145 => X"9F43",
	146 => X"9656",
	147 => X"8ECA",
	148 => X"88B8",
	149 => X"8434",
	150 => X"814D",
	151 => X"800D",
	152 => X"8078",
	153 => X"828C",
	154 => X"8643",
	155 => X"8B91",
	156 => X"9263",
	157 => X"9AA2",
	158 => X"A434",
	159 => X"AEF9",
	160 => X"BACB",
	161 => X"C785",
	162 => X"D4FB",
	163 => X"E301",
	164 => X"F167",
	165 => X"FFFE",
	166 => X"0E97",
	167 => X"1CFD",
	168 => X"2B03",
	169 => X"3879",
	170 => X"4533",
	171 => X"5105",
	172 => X"5BCA",
	173 => X"655C",
	174 => X"6D9B",
	175 => X"746D",
	176 => X"79BB",
	177 => X"7D72",
	178 => X"7F86",
	179 => X"7FF1",
	180 => X"7EB1",
	181 => X"7BCA",
	182 => X"7746",
	183 => X"7134",
	184 => X"69A8",
	185 => X"60BB",
	186 => X"568C",
	187 => X"4B3B",
	188 => X"3EF0",
	189 => X"31D3",
	190 => X"240F",
	191 => X"15D3",
	192 => X"074E",
	193 => X"F8B0",
	194 => X"EA2B",
	195 => X"DBEF",
	196 => X"CE2B",
	197 => X"C10E",
	198 => X"B4C3",
	199 => X"A972",
	200 => X"9F43",
	201 => X"9656",
	202 => X"8ECA",
	203 => X"88B8",
	204 => X"8434",
	205 => X"814D",
	206 => X"800D",
	207 => X"8078",
	208 => X"828C",
	209 => X"8643",
	210 => X"8B91",
	211 => X"9263",
	212 => X"9AA2",
	213 => X"A434",
	214 => X"AEF9",
	215 => X"BACB",
	216 => X"C785",
	217 => X"D4FB",
	218 => X"E301",
	219 => X"F167",
	220 => X"FFFE",
	221 => X"0E97",
	222 => X"1CFD",
	223 => X"2B03",
	224 => X"3879",
	225 => X"4533",
	226 => X"5105",
	227 => X"5BCA",
	228 => X"655C",
	229 => X"6D9B",
	230 => X"746D",
	231 => X"79BB",
	232 => X"7D72",
	233 => X"7F86",
	234 => X"7FF1",
	235 => X"7EB1",
	236 => X"7BCA",
	237 => X"7746",
	238 => X"7134",
	239 => X"69A8",
	240 => X"60BB",
	241 => X"568C",
	242 => X"4B3B",
	243 => X"3EF0",
	244 => X"31D3",
	245 => X"240F",
	246 => X"15D3",
	247 => X"074E",
	others => X"0000"
);

CONSTANT DS5: hex := (
	000 => X"0000",
	001 => X"0F6D",
	002 => X"1EA1",
	003 => X"2D63",
	004 => X"3B7B",
	005 => X"48B5",
	006 => X"54E0",
	007 => X"5FCE",
	008 => X"6956",
	009 => X"7155",
	010 => X"77AD",
	011 => X"7C46",
	012 => X"7F10",
	013 => X"7FFF",
	014 => X"7F10",
	015 => X"7C46",
	016 => X"77AD",
	017 => X"7155",
	018 => X"6956",
	019 => X"5FCE",
	020 => X"54E0",
	021 => X"48B5",
	022 => X"3B7B",
	023 => X"2D63",
	024 => X"1EA1",
	025 => X"0F6D",
	026 => X"FFFE",
	027 => X"F091",
	028 => X"E15D",
	029 => X"D29B",
	030 => X"C483",
	031 => X"B749",
	032 => X"AB1E",
	033 => X"A030",
	034 => X"96A8",
	035 => X"8EA9",
	036 => X"8851",
	037 => X"83B8",
	038 => X"80EE",
	039 => X"8000",
	040 => X"80EE",
	041 => X"83B8",
	042 => X"8851",
	043 => X"8EA9",
	044 => X"96A8",
	045 => X"A030",
	046 => X"AB1E",
	047 => X"B749",
	048 => X"C483",
	049 => X"D29B",
	050 => X"E15D",
	051 => X"F091",
	052 => X"FFFE",
	053 => X"0F6D",
	054 => X"1EA1",
	055 => X"2D63",
	056 => X"3B7B",
	057 => X"48B5",
	058 => X"54E0",
	059 => X"5FCE",
	060 => X"6956",
	061 => X"7155",
	062 => X"77AD",
	063 => X"7C46",
	064 => X"7F10",
	065 => X"7FFF",
	066 => X"7F10",
	067 => X"7C46",
	068 => X"77AD",
	069 => X"7155",
	070 => X"6956",
	071 => X"5FCE",
	072 => X"54E0",
	073 => X"48B5",
	074 => X"3B7B",
	075 => X"2D63",
	076 => X"1EA1",
	077 => X"0F6D",
	078 => X"0000",
	079 => X"F091",
	080 => X"E15D",
	081 => X"D29B",
	082 => X"C483",
	083 => X"B749",
	084 => X"AB1E",
	085 => X"A030",
	086 => X"96A8",
	087 => X"8EA9",
	088 => X"8851",
	089 => X"83B8",
	090 => X"80EE",
	091 => X"8000",
	092 => X"80EE",
	093 => X"83B8",
	094 => X"8851",
	095 => X"8EA9",
	096 => X"96A8",
	097 => X"A030",
	098 => X"AB1E",
	099 => X"B749",
	100 => X"C483",
	101 => X"D29B",
	102 => X"E15D",
	103 => X"F091",
	104 => X"FFFE",
	105 => X"0F6D",
	106 => X"1EA1",
	107 => X"2D63",
	108 => X"3B7B",
	109 => X"48B5",
	110 => X"54E0",
	111 => X"5FCE",
	112 => X"6956",
	113 => X"7155",
	114 => X"77AD",
	115 => X"7C46",
	116 => X"7F10",
	117 => X"7FFF",
	118 => X"7F10",
	119 => X"7C46",
	120 => X"77AD",
	121 => X"7155",
	122 => X"6956",
	123 => X"5FCE",
	124 => X"54E0",
	125 => X"48B5",
	126 => X"3B7B",
	127 => X"2D63",
	128 => X"1EA1",
	129 => X"0F6D",
	130 => X"0000",
	131 => X"F091",
	132 => X"E15D",
	133 => X"D29B",
	134 => X"C483",
	135 => X"B749",
	136 => X"AB1E",
	137 => X"A030",
	138 => X"96A8",
	139 => X"8EA9",
	140 => X"8851",
	141 => X"83B8",
	142 => X"80EE",
	143 => X"8000",
	144 => X"80EE",
	145 => X"83B8",
	146 => X"8851",
	147 => X"8EA9",
	148 => X"96A8",
	149 => X"A030",
	150 => X"AB1E",
	151 => X"B749",
	152 => X"C483",
	153 => X"D29B",
	154 => X"E15D",
	155 => X"F091",
	156 => X"FFFE",
	157 => X"0F6D",
	158 => X"1EA1",
	159 => X"2D63",
	160 => X"3B7B",
	161 => X"48B5",
	162 => X"54E0",
	163 => X"5FCE",
	164 => X"6956",
	165 => X"7155",
	166 => X"77AD",
	167 => X"7C46",
	168 => X"7F10",
	169 => X"7FFF",
	170 => X"7F10",
	171 => X"7C46",
	172 => X"77AD",
	173 => X"7155",
	174 => X"6956",
	175 => X"5FCE",
	176 => X"54E0",
	177 => X"48B5",
	178 => X"3B7B",
	179 => X"2D63",
	180 => X"1EA1",
	181 => X"0F6D",
	182 => X"0000",
	183 => X"F091",
	184 => X"E15D",
	185 => X"D29B",
	186 => X"C483",
	187 => X"B749",
	188 => X"AB1E",
	189 => X"A030",
	190 => X"96A8",
	191 => X"8EA9",
	192 => X"8851",
	193 => X"83B8",
	194 => X"80EE",
	195 => X"8000",
	196 => X"80EE",
	197 => X"83B8",
	198 => X"8851",
	199 => X"8EA9",
	200 => X"96A8",
	201 => X"A030",
	202 => X"AB1E",
	203 => X"B749",
	204 => X"C483",
	205 => X"D29B",
	206 => X"E15D",
	207 => X"F091",
	208 => X"FFFE",
	209 => X"0F6D",
	210 => X"1EA1",
	211 => X"2D63",
	212 => X"3B7B",
	213 => X"48B5",
	214 => X"54E0",
	215 => X"5FCE",
	216 => X"6956",
	217 => X"7155",
	218 => X"77AD",
	219 => X"7C46",
	220 => X"7F10",
	221 => X"7FFF",
	222 => X"7F10",
	223 => X"7C46",
	224 => X"77AD",
	225 => X"7155",
	226 => X"6956",
	227 => X"5FCE",
	228 => X"54E0",
	229 => X"48B5",
	230 => X"3B7B",
	231 => X"2D63",
	232 => X"1EA1",
	233 => X"0F6D",
	234 => X"0000",
	235 => X"F091",
	236 => X"E15D",
	237 => X"D29B",
	238 => X"C483",
	239 => X"B749",
	240 => X"AB1E",
	241 => X"A030",
	242 => X"96A8",
	243 => X"8EA9",
	244 => X"8851",
	245 => X"83B8",
	246 => X"80EE",
	247 => X"8000",
	others => X"0000"
);

CONSTANT E5: hex := (
	000 => X"0000",
	001 => X"105E",
	002 => X"2077",
	003 => X"3008",
	004 => X"3ECF",
	005 => X"4C8E",
	006 => X"590B",
	007 => X"6412",
	008 => X"6D74",
	009 => X"750A",
	010 => X"7AB4",
	011 => X"7E5A",
	012 => X"7FEE",
	013 => X"7F67",
	014 => X"7CC9",
	015 => X"781E",
	016 => X"717B",
	017 => X"68FA",
	018 => X"5EC0",
	019 => X"52F8",
	020 => X"45D3",
	021 => X"3789",
	022 => X"2855",
	023 => X"1877",
	024 => X"0833",
	025 => X"F7CB",
	026 => X"E787",
	027 => X"D7A9",
	028 => X"C875",
	029 => X"BA2B",
	030 => X"AD06",
	031 => X"A13E",
	032 => X"9704",
	033 => X"8E83",
	034 => X"87E0",
	035 => X"8335",
	036 => X"8097",
	037 => X"8010",
	038 => X"81A4",
	039 => X"854A",
	040 => X"8AF4",
	041 => X"928A",
	042 => X"9BEC",
	043 => X"A6F3",
	044 => X"B370",
	045 => X"C12F",
	046 => X"CFF6",
	047 => X"DF87",
	048 => X"EFA0",
	049 => X"FFFE",
	050 => X"105E",
	051 => X"2077",
	052 => X"3008",
	053 => X"3ECF",
	054 => X"4C8E",
	055 => X"590B",
	056 => X"6412",
	057 => X"6D74",
	058 => X"750A",
	059 => X"7AB4",
	060 => X"7E5A",
	061 => X"7FEE",
	062 => X"7F67",
	063 => X"7CC9",
	064 => X"781E",
	065 => X"717B",
	066 => X"68FA",
	067 => X"5EC0",
	068 => X"52F8",
	069 => X"45D3",
	070 => X"3789",
	071 => X"2855",
	072 => X"1877",
	073 => X"0833",
	074 => X"F7CB",
	075 => X"E787",
	076 => X"D7A9",
	077 => X"C875",
	078 => X"BA2B",
	079 => X"AD06",
	080 => X"A13E",
	081 => X"9704",
	082 => X"8E83",
	083 => X"87E0",
	084 => X"8335",
	085 => X"8097",
	086 => X"8010",
	087 => X"81A4",
	088 => X"854A",
	089 => X"8AF4",
	090 => X"928A",
	091 => X"9BEC",
	092 => X"A6F3",
	093 => X"B370",
	094 => X"C12F",
	095 => X"CFF6",
	096 => X"DF87",
	097 => X"EFA0",
	098 => X"0000",
	099 => X"105E",
	100 => X"2077",
	101 => X"3008",
	102 => X"3ECF",
	103 => X"4C8E",
	104 => X"590B",
	105 => X"6412",
	106 => X"6D74",
	107 => X"750A",
	108 => X"7AB4",
	109 => X"7E5A",
	110 => X"7FEE",
	111 => X"7F67",
	112 => X"7CC9",
	113 => X"781E",
	114 => X"717B",
	115 => X"68FA",
	116 => X"5EC0",
	117 => X"52F8",
	118 => X"45D3",
	119 => X"3789",
	120 => X"2855",
	121 => X"1877",
	122 => X"0833",
	123 => X"F7CB",
	124 => X"E787",
	125 => X"D7A9",
	126 => X"C875",
	127 => X"BA2B",
	128 => X"AD06",
	129 => X"A13E",
	130 => X"9704",
	131 => X"8E83",
	132 => X"87E0",
	133 => X"8335",
	134 => X"8097",
	135 => X"8010",
	136 => X"81A4",
	137 => X"854A",
	138 => X"8AF4",
	139 => X"928A",
	140 => X"9BEC",
	141 => X"A6F3",
	142 => X"B370",
	143 => X"C12F",
	144 => X"CFF6",
	145 => X"DF87",
	146 => X"EFA0",
	147 => X"0000",
	148 => X"105E",
	149 => X"2077",
	150 => X"3008",
	151 => X"3ECF",
	152 => X"4C8E",
	153 => X"590B",
	154 => X"6412",
	155 => X"6D74",
	156 => X"750A",
	157 => X"7AB4",
	158 => X"7E5A",
	159 => X"7FEE",
	160 => X"7F67",
	161 => X"7CC9",
	162 => X"781E",
	163 => X"717B",
	164 => X"68FA",
	165 => X"5EC0",
	166 => X"52F8",
	167 => X"45D3",
	168 => X"3789",
	169 => X"2855",
	170 => X"1877",
	171 => X"0833",
	172 => X"F7CB",
	173 => X"E787",
	174 => X"D7A9",
	175 => X"C875",
	176 => X"BA2B",
	177 => X"AD06",
	178 => X"A13E",
	179 => X"9704",
	180 => X"8E83",
	181 => X"87E0",
	182 => X"8335",
	183 => X"8097",
	184 => X"8010",
	185 => X"81A4",
	186 => X"854A",
	187 => X"8AF4",
	188 => X"928A",
	189 => X"9BEC",
	190 => X"A6F3",
	191 => X"B370",
	192 => X"C12F",
	193 => X"CFF6",
	194 => X"DF87",
	195 => X"EFA0",
	196 => X"FFFE",
	197 => X"105E",
	198 => X"2077",
	199 => X"3008",
	200 => X"3ECF",
	201 => X"4C8E",
	202 => X"590B",
	203 => X"6412",
	204 => X"6D74",
	205 => X"750A",
	206 => X"7AB4",
	207 => X"7E5A",
	208 => X"7FEE",
	209 => X"7F67",
	210 => X"7CC9",
	211 => X"781E",
	212 => X"717B",
	213 => X"68FA",
	214 => X"5EC0",
	215 => X"52F8",
	216 => X"45D3",
	217 => X"3789",
	218 => X"2855",
	219 => X"1877",
	220 => X"0833",
	221 => X"F7CB",
	222 => X"E787",
	223 => X"D7A9",
	224 => X"C875",
	225 => X"BA2B",
	226 => X"AD06",
	227 => X"A13E",
	228 => X"9704",
	229 => X"8E83",
	230 => X"87E0",
	231 => X"8335",
	232 => X"8097",
	233 => X"8010",
	234 => X"81A4",
	235 => X"854A",
	236 => X"8AF4",
	237 => X"928A",
	238 => X"9BEC",
	239 => X"A6F3",
	240 => X"B370",
	241 => X"C12F",
	242 => X"CFF6",
	243 => X"DF87",
	244 => X"EFA0",
	245 => X"FFFE",
	246 => X"105E",
	247 => X"2077",
	others => X"0000"
);

CONSTANT F5: hex := (
	000 => X"0000",
	001 => X"110F",
	002 => X"21D0",
	003 => X"31F7",
	004 => X"413A",
	005 => X"4F53",
	006 => X"5C01",
	007 => X"670B",
	008 => X"703F",
	009 => X"7771",
	010 => X"7C82",
	011 => X"7F5A",
	012 => X"7FEC",
	013 => X"7E36",
	014 => X"7A3F",
	015 => X"741A",
	016 => X"6BE3",
	017 => X"61BE",
	018 => X"55DB",
	019 => X"4870",
	020 => X"39BA",
	021 => X"29FC",
	022 => X"197E",
	023 => X"088C",
	024 => X"F772",
	025 => X"E680",
	026 => X"D602",
	027 => X"C644",
	028 => X"B78E",
	029 => X"AA23",
	030 => X"9E40",
	031 => X"941B",
	032 => X"8BE4",
	033 => X"85BF",
	034 => X"81C8",
	035 => X"8012",
	036 => X"80A4",
	037 => X"837C",
	038 => X"888D",
	039 => X"8FBF",
	040 => X"98F3",
	041 => X"A3FD",
	042 => X"B0AB",
	043 => X"BEC4",
	044 => X"CE07",
	045 => X"DE2E",
	046 => X"EEEF",
	047 => X"0000",
	048 => X"110F",
	049 => X"21D0",
	050 => X"31F7",
	051 => X"413A",
	052 => X"4F53",
	053 => X"5C01",
	054 => X"670B",
	055 => X"703F",
	056 => X"7771",
	057 => X"7C82",
	058 => X"7F5A",
	059 => X"7FEC",
	060 => X"7E36",
	061 => X"7A3F",
	062 => X"741A",
	063 => X"6BE3",
	064 => X"61BE",
	065 => X"55DB",
	066 => X"4870",
	067 => X"39BA",
	068 => X"29FC",
	069 => X"197E",
	070 => X"088C",
	071 => X"F772",
	072 => X"E680",
	073 => X"D602",
	074 => X"C644",
	075 => X"B78E",
	076 => X"AA23",
	077 => X"9E40",
	078 => X"941B",
	079 => X"8BE4",
	080 => X"85BF",
	081 => X"81C8",
	082 => X"8012",
	083 => X"80A4",
	084 => X"837C",
	085 => X"888D",
	086 => X"8FBF",
	087 => X"98F3",
	088 => X"A3FD",
	089 => X"B0AB",
	090 => X"BEC4",
	091 => X"CE07",
	092 => X"DE2E",
	093 => X"EEEF",
	094 => X"0000",
	095 => X"110F",
	096 => X"21D0",
	097 => X"31F7",
	098 => X"413A",
	099 => X"4F53",
	100 => X"5C01",
	101 => X"670B",
	102 => X"703F",
	103 => X"7771",
	104 => X"7C82",
	105 => X"7F5A",
	106 => X"7FEC",
	107 => X"7E36",
	108 => X"7A3F",
	109 => X"741A",
	110 => X"6BE3",
	111 => X"61BE",
	112 => X"55DB",
	113 => X"4870",
	114 => X"39BA",
	115 => X"29FC",
	116 => X"197E",
	117 => X"088C",
	118 => X"F772",
	119 => X"E680",
	120 => X"D602",
	121 => X"C644",
	122 => X"B78E",
	123 => X"AA23",
	124 => X"9E40",
	125 => X"941B",
	126 => X"8BE4",
	127 => X"85BF",
	128 => X"81C8",
	129 => X"8012",
	130 => X"80A4",
	131 => X"837C",
	132 => X"888D",
	133 => X"8FBF",
	134 => X"98F3",
	135 => X"A3FD",
	136 => X"B0AB",
	137 => X"BEC4",
	138 => X"CE07",
	139 => X"DE2E",
	140 => X"EEEF",
	141 => X"0000",
	142 => X"110F",
	143 => X"21D0",
	144 => X"31F7",
	145 => X"413A",
	146 => X"4F53",
	147 => X"5C01",
	148 => X"670B",
	149 => X"703F",
	150 => X"7771",
	151 => X"7C82",
	152 => X"7F5A",
	153 => X"7FEC",
	154 => X"7E36",
	155 => X"7A3F",
	156 => X"741A",
	157 => X"6BE3",
	158 => X"61BE",
	159 => X"55DB",
	160 => X"4870",
	161 => X"39BA",
	162 => X"29FC",
	163 => X"197E",
	164 => X"088C",
	165 => X"F772",
	166 => X"E680",
	167 => X"D602",
	168 => X"C644",
	169 => X"B78E",
	170 => X"AA23",
	171 => X"9E40",
	172 => X"941B",
	173 => X"8BE4",
	174 => X"85BF",
	175 => X"81C8",
	176 => X"8012",
	177 => X"80A4",
	178 => X"837C",
	179 => X"888D",
	180 => X"8FBF",
	181 => X"98F3",
	182 => X"A3FD",
	183 => X"B0AB",
	184 => X"BEC4",
	185 => X"CE07",
	186 => X"DE2E",
	187 => X"EEEF",
	188 => X"0000",
	189 => X"110F",
	190 => X"21D0",
	191 => X"31F7",
	192 => X"413A",
	193 => X"4F53",
	194 => X"5C01",
	195 => X"670B",
	196 => X"703F",
	197 => X"7771",
	198 => X"7C82",
	199 => X"7F5A",
	200 => X"7FEC",
	201 => X"7E36",
	202 => X"7A3F",
	203 => X"741A",
	204 => X"6BE3",
	205 => X"61BE",
	206 => X"55DB",
	207 => X"4870",
	208 => X"39BA",
	209 => X"29FC",
	210 => X"197E",
	211 => X"088C",
	212 => X"F772",
	213 => X"E680",
	214 => X"D602",
	215 => X"C644",
	216 => X"B78E",
	217 => X"AA23",
	218 => X"9E40",
	219 => X"941B",
	220 => X"8BE4",
	221 => X"85BF",
	222 => X"81C8",
	223 => X"8012",
	224 => X"80A4",
	225 => X"837C",
	226 => X"888D",
	227 => X"8FBF",
	228 => X"98F3",
	229 => X"A3FD",
	230 => X"B0AB",
	231 => X"BEC4",
	232 => X"CE07",
	233 => X"DE2E",
	234 => X"EEEF",
	235 => X"0000",
	236 => X"110F",
	237 => X"21D0",
	238 => X"31F7",
	239 => X"413A",
	240 => X"4F53",
	241 => X"5C01",
	242 => X"670B",
	243 => X"703F",
	244 => X"7771",
	245 => X"7C82",
	246 => X"7F5A",
	247 => X"7FEC",
	others => X"0000"
);

CONSTANT FS5: hex := (
	000 => X"0000",
	001 => X"1237",
	002 => X"240F",
	003 => X"352B",
	004 => X"4533",
	005 => X"53D1",
	006 => X"60BB",
	007 => X"6BAD",
	008 => X"746D",
	009 => X"7ACF",
	010 => X"7EB1",
	011 => X"7FFF",
	012 => X"7EB1",
	013 => X"7ACF",
	014 => X"746D",
	015 => X"6BAD",
	016 => X"60BB",
	017 => X"53D1",
	018 => X"4533",
	019 => X"352B",
	020 => X"240F",
	021 => X"1237",
	022 => X"FFFE",
	023 => X"EDC7",
	024 => X"DBEF",
	025 => X"CAD3",
	026 => X"BACB",
	027 => X"AC2D",
	028 => X"9F43",
	029 => X"9451",
	030 => X"8B91",
	031 => X"852F",
	032 => X"814D",
	033 => X"8000",
	034 => X"814D",
	035 => X"852F",
	036 => X"8B91",
	037 => X"9451",
	038 => X"9F43",
	039 => X"AC2D",
	040 => X"BACB",
	041 => X"CAD3",
	042 => X"DBEF",
	043 => X"EDC7",
	044 => X"0000",
	045 => X"1237",
	046 => X"240F",
	047 => X"352B",
	048 => X"4533",
	049 => X"53D1",
	050 => X"60BB",
	051 => X"6BAD",
	052 => X"746D",
	053 => X"7ACF",
	054 => X"7EB1",
	055 => X"7FFF",
	056 => X"7EB1",
	057 => X"7ACF",
	058 => X"746D",
	059 => X"6BAD",
	060 => X"60BB",
	061 => X"53D1",
	062 => X"4533",
	063 => X"352B",
	064 => X"240F",
	065 => X"1237",
	066 => X"FFFE",
	067 => X"EDC7",
	068 => X"DBEF",
	069 => X"CAD3",
	070 => X"BACB",
	071 => X"AC2D",
	072 => X"9F43",
	073 => X"9451",
	074 => X"8B91",
	075 => X"852F",
	076 => X"814D",
	077 => X"8000",
	078 => X"814D",
	079 => X"852F",
	080 => X"8B91",
	081 => X"9451",
	082 => X"9F43",
	083 => X"AC2D",
	084 => X"BACB",
	085 => X"CAD3",
	086 => X"DBEF",
	087 => X"EDC7",
	088 => X"FFFE",
	089 => X"1237",
	090 => X"240F",
	091 => X"352B",
	092 => X"4533",
	093 => X"53D1",
	094 => X"60BB",
	095 => X"6BAD",
	096 => X"746D",
	097 => X"7ACF",
	098 => X"7EB1",
	099 => X"7FFF",
	100 => X"7EB1",
	101 => X"7ACF",
	102 => X"746D",
	103 => X"6BAD",
	104 => X"60BB",
	105 => X"53D1",
	106 => X"4533",
	107 => X"352B",
	108 => X"240F",
	109 => X"1237",
	110 => X"0000",
	111 => X"EDC7",
	112 => X"DBEF",
	113 => X"CAD3",
	114 => X"BACB",
	115 => X"AC2D",
	116 => X"9F43",
	117 => X"9451",
	118 => X"8B91",
	119 => X"852F",
	120 => X"814D",
	121 => X"8000",
	122 => X"814D",
	123 => X"852F",
	124 => X"8B91",
	125 => X"9451",
	126 => X"9F43",
	127 => X"AC2D",
	128 => X"BACB",
	129 => X"CAD3",
	130 => X"DBEF",
	131 => X"EDC7",
	132 => X"FFFE",
	133 => X"1237",
	134 => X"240F",
	135 => X"352B",
	136 => X"4533",
	137 => X"53D1",
	138 => X"60BB",
	139 => X"6BAD",
	140 => X"746D",
	141 => X"7ACF",
	142 => X"7EB1",
	143 => X"7FFF",
	144 => X"7EB1",
	145 => X"7ACF",
	146 => X"746D",
	147 => X"6BAD",
	148 => X"60BB",
	149 => X"53D1",
	150 => X"4533",
	151 => X"352B",
	152 => X"240F",
	153 => X"1237",
	154 => X"0000",
	155 => X"EDC7",
	156 => X"DBEF",
	157 => X"CAD3",
	158 => X"BACB",
	159 => X"AC2D",
	160 => X"9F43",
	161 => X"9451",
	162 => X"8B91",
	163 => X"852F",
	164 => X"814D",
	165 => X"8000",
	166 => X"814D",
	167 => X"852F",
	168 => X"8B91",
	169 => X"9451",
	170 => X"9F43",
	171 => X"AC2D",
	172 => X"BACB",
	173 => X"CAD3",
	174 => X"DBEF",
	175 => X"EDC7",
	176 => X"0000",
	177 => X"1237",
	178 => X"240F",
	179 => X"352B",
	180 => X"4533",
	181 => X"53D1",
	182 => X"60BB",
	183 => X"6BAD",
	184 => X"746D",
	185 => X"7ACF",
	186 => X"7EB1",
	187 => X"7FFF",
	188 => X"7EB1",
	189 => X"7ACF",
	190 => X"746D",
	191 => X"6BAD",
	192 => X"60BB",
	193 => X"53D1",
	194 => X"4533",
	195 => X"352B",
	196 => X"240F",
	197 => X"1237",
	198 => X"FFFE",
	199 => X"EDC7",
	200 => X"DBEF",
	201 => X"CAD3",
	202 => X"BACB",
	203 => X"AC2D",
	204 => X"9F43",
	205 => X"9451",
	206 => X"8B91",
	207 => X"852F",
	208 => X"814D",
	209 => X"8000",
	210 => X"814D",
	211 => X"852F",
	212 => X"8B91",
	213 => X"9451",
	214 => X"9F43",
	215 => X"AC2D",
	216 => X"BACB",
	217 => X"CAD3",
	218 => X"DBEF",
	219 => X"EDC7",
	220 => X"0000",
	221 => X"1237",
	222 => X"240F",
	223 => X"352B",
	224 => X"4533",
	225 => X"53D1",
	226 => X"60BB",
	227 => X"6BAD",
	228 => X"746D",
	229 => X"7ACF",
	230 => X"7EB1",
	231 => X"7FFF",
	232 => X"7EB1",
	233 => X"7ACF",
	234 => X"746D",
	235 => X"6BAD",
	236 => X"60BB",
	237 => X"53D1",
	238 => X"4533",
	239 => X"352B",
	240 => X"240F",
	241 => X"1237",
	242 => X"FFFE",
	243 => X"EDC7",
	244 => X"DBEF",
	245 => X"CAD3",
	246 => X"BACB",
	247 => X"AC2D",
	others => X"0000"
);

CONSTANT G5: hex := (
	000 => X"0000",
	001 => X"1313",
	002 => X"25BA",
	003 => X"3789",
	004 => X"481A",
	005 => X"570F",
	006 => X"6412",
	007 => X"6ED9",
	008 => X"7725",
	009 => X"7CC9",
	010 => X"7FA3",
	011 => X"7FA3",
	012 => X"7CC9",
	013 => X"7725",
	014 => X"6ED9",
	015 => X"6412",
	016 => X"570F",
	017 => X"481A",
	018 => X"3789",
	019 => X"25BA",
	020 => X"1313",
	021 => X"FFFE",
	022 => X"ECEB",
	023 => X"DA44",
	024 => X"C875",
	025 => X"B7E4",
	026 => X"A8EF",
	027 => X"9BEC",
	028 => X"9125",
	029 => X"88D9",
	030 => X"8335",
	031 => X"805B",
	032 => X"805B",
	033 => X"8335",
	034 => X"88D9",
	035 => X"9125",
	036 => X"9BEC",
	037 => X"A8EF",
	038 => X"B7E4",
	039 => X"C875",
	040 => X"DA44",
	041 => X"ECEB",
	042 => X"FFFE",
	043 => X"1313",
	044 => X"25BA",
	045 => X"3789",
	046 => X"481A",
	047 => X"570F",
	048 => X"6412",
	049 => X"6ED9",
	050 => X"7725",
	051 => X"7CC9",
	052 => X"7FA3",
	053 => X"7FA3",
	054 => X"7CC9",
	055 => X"7725",
	056 => X"6ED9",
	057 => X"6412",
	058 => X"570F",
	059 => X"481A",
	060 => X"3789",
	061 => X"25BA",
	062 => X"1313",
	063 => X"0000",
	064 => X"ECEB",
	065 => X"DA44",
	066 => X"C875",
	067 => X"B7E4",
	068 => X"A8EF",
	069 => X"9BEC",
	070 => X"9125",
	071 => X"88D9",
	072 => X"8335",
	073 => X"805B",
	074 => X"805B",
	075 => X"8335",
	076 => X"88D9",
	077 => X"9125",
	078 => X"9BEC",
	079 => X"A8EF",
	080 => X"B7E4",
	081 => X"C875",
	082 => X"DA44",
	083 => X"ECEB",
	084 => X"FFFE",
	085 => X"1313",
	086 => X"25BA",
	087 => X"3789",
	088 => X"481A",
	089 => X"570F",
	090 => X"6412",
	091 => X"6ED9",
	092 => X"7725",
	093 => X"7CC9",
	094 => X"7FA3",
	095 => X"7FA3",
	096 => X"7CC9",
	097 => X"7725",
	098 => X"6ED9",
	099 => X"6412",
	100 => X"570F",
	101 => X"481A",
	102 => X"3789",
	103 => X"25BA",
	104 => X"1313",
	105 => X"0000",
	106 => X"ECEB",
	107 => X"DA44",
	108 => X"C875",
	109 => X"B7E4",
	110 => X"A8EF",
	111 => X"9BEC",
	112 => X"9125",
	113 => X"88D9",
	114 => X"8335",
	115 => X"805B",
	116 => X"805B",
	117 => X"8335",
	118 => X"88D9",
	119 => X"9125",
	120 => X"9BEC",
	121 => X"A8EF",
	122 => X"B7E4",
	123 => X"C875",
	124 => X"DA44",
	125 => X"ECEB",
	126 => X"FFFE",
	127 => X"1313",
	128 => X"25BA",
	129 => X"3789",
	130 => X"481A",
	131 => X"570F",
	132 => X"6412",
	133 => X"6ED9",
	134 => X"7725",
	135 => X"7CC9",
	136 => X"7FA3",
	137 => X"7FA3",
	138 => X"7CC9",
	139 => X"7725",
	140 => X"6ED9",
	141 => X"6412",
	142 => X"570F",
	143 => X"481A",
	144 => X"3789",
	145 => X"25BA",
	146 => X"1313",
	147 => X"FFFE",
	148 => X"ECEB",
	149 => X"DA44",
	150 => X"C875",
	151 => X"B7E4",
	152 => X"A8EF",
	153 => X"9BEC",
	154 => X"9125",
	155 => X"88D9",
	156 => X"8335",
	157 => X"805B",
	158 => X"805B",
	159 => X"8335",
	160 => X"88D9",
	161 => X"9125",
	162 => X"9BEC",
	163 => X"A8EF",
	164 => X"B7E4",
	165 => X"C875",
	166 => X"DA44",
	167 => X"ECEB",
	168 => X"0000",
	169 => X"1313",
	170 => X"25BA",
	171 => X"3789",
	172 => X"481A",
	173 => X"570F",
	174 => X"6412",
	175 => X"6ED9",
	176 => X"7725",
	177 => X"7CC9",
	178 => X"7FA3",
	179 => X"7FA3",
	180 => X"7CC9",
	181 => X"7725",
	182 => X"6ED9",
	183 => X"6412",
	184 => X"570F",
	185 => X"481A",
	186 => X"3789",
	187 => X"25BA",
	188 => X"1313",
	189 => X"FFFE",
	190 => X"ECEB",
	191 => X"DA44",
	192 => X"C875",
	193 => X"B7E4",
	194 => X"A8EF",
	195 => X"9BEC",
	196 => X"9125",
	197 => X"88D9",
	198 => X"8335",
	199 => X"805B",
	200 => X"805B",
	201 => X"8335",
	202 => X"88D9",
	203 => X"9125",
	204 => X"9BEC",
	205 => X"A8EF",
	206 => X"B7E4",
	207 => X"C875",
	208 => X"DA44",
	209 => X"ECEB",
	210 => X"0000",
	211 => X"1313",
	212 => X"25BA",
	213 => X"3789",
	214 => X"481A",
	215 => X"570F",
	216 => X"6412",
	217 => X"6ED9",
	218 => X"7725",
	219 => X"7CC9",
	220 => X"7FA3",
	221 => X"7FA3",
	222 => X"7CC9",
	223 => X"7725",
	224 => X"6ED9",
	225 => X"6412",
	226 => X"570F",
	227 => X"481A",
	228 => X"3789",
	229 => X"25BA",
	230 => X"1313",
	231 => X"FFFE",
	232 => X"ECEB",
	233 => X"DA44",
	234 => X"C875",
	235 => X"B7E4",
	236 => X"A8EF",
	237 => X"9BEC",
	238 => X"9125",
	239 => X"88D9",
	240 => X"8335",
	241 => X"805B",
	242 => X"805B",
	243 => X"8335",
	244 => X"88D9",
	245 => X"9125",
	246 => X"9BEC",
	247 => X"A8EF",
	others => X"0000"
);

CONSTANT GS5: hex := (
	000 => X"0000",
	001 => X"1488",
	002 => X"2888",
	003 => X"3B7B",
	004 => X"4CE4",
	005 => X"5C4F",
	006 => X"6956",
	007 => X"73A3",
	008 => X"7AF1",
	009 => X"7F10",
	010 => X"7FE4",
	011 => X"7D68",
	012 => X"77AD",
	013 => X"6ED9",
	014 => X"6325",
	015 => X"54E0",
	016 => X"4468",
	017 => X"322B",
	018 => X"1EA1",
	019 => X"0A4C",
	020 => X"F5B2",
	021 => X"E15D",
	022 => X"CDD3",
	023 => X"BB96",
	024 => X"AB1E",
	025 => X"9CD9",
	026 => X"9125",
	027 => X"8851",
	028 => X"8296",
	029 => X"801A",
	030 => X"80EE",
	031 => X"850D",
	032 => X"8C5B",
	033 => X"96A8",
	034 => X"A3AF",
	035 => X"B31A",
	036 => X"C483",
	037 => X"D776",
	038 => X"EB76",
	039 => X"FFFE",
	040 => X"1488",
	041 => X"2888",
	042 => X"3B7B",
	043 => X"4CE4",
	044 => X"5C4F",
	045 => X"6956",
	046 => X"73A3",
	047 => X"7AF1",
	048 => X"7F10",
	049 => X"7FE4",
	050 => X"7D68",
	051 => X"77AD",
	052 => X"6ED9",
	053 => X"6325",
	054 => X"54E0",
	055 => X"4468",
	056 => X"322B",
	057 => X"1EA1",
	058 => X"0A4C",
	059 => X"F5B2",
	060 => X"E15D",
	061 => X"CDD3",
	062 => X"BB96",
	063 => X"AB1E",
	064 => X"9CD9",
	065 => X"9125",
	066 => X"8851",
	067 => X"8296",
	068 => X"801A",
	069 => X"80EE",
	070 => X"850D",
	071 => X"8C5B",
	072 => X"96A8",
	073 => X"A3AF",
	074 => X"B31A",
	075 => X"C483",
	076 => X"D776",
	077 => X"EB76",
	078 => X"0000",
	079 => X"1488",
	080 => X"2888",
	081 => X"3B7B",
	082 => X"4CE4",
	083 => X"5C4F",
	084 => X"6956",
	085 => X"73A3",
	086 => X"7AF1",
	087 => X"7F10",
	088 => X"7FE4",
	089 => X"7D68",
	090 => X"77AD",
	091 => X"6ED9",
	092 => X"6325",
	093 => X"54E0",
	094 => X"4468",
	095 => X"322B",
	096 => X"1EA1",
	097 => X"0A4C",
	098 => X"F5B2",
	099 => X"E15D",
	100 => X"CDD3",
	101 => X"BB96",
	102 => X"AB1E",
	103 => X"9CD9",
	104 => X"9125",
	105 => X"8851",
	106 => X"8296",
	107 => X"801A",
	108 => X"80EE",
	109 => X"850D",
	110 => X"8C5B",
	111 => X"96A8",
	112 => X"A3AF",
	113 => X"B31A",
	114 => X"C483",
	115 => X"D776",
	116 => X"EB76",
	117 => X"0000",
	118 => X"1488",
	119 => X"2888",
	120 => X"3B7B",
	121 => X"4CE4",
	122 => X"5C4F",
	123 => X"6956",
	124 => X"73A3",
	125 => X"7AF1",
	126 => X"7F10",
	127 => X"7FE4",
	128 => X"7D68",
	129 => X"77AD",
	130 => X"6ED9",
	131 => X"6325",
	132 => X"54E0",
	133 => X"4468",
	134 => X"322B",
	135 => X"1EA1",
	136 => X"0A4C",
	137 => X"F5B2",
	138 => X"E15D",
	139 => X"CDD3",
	140 => X"BB96",
	141 => X"AB1E",
	142 => X"9CD9",
	143 => X"9125",
	144 => X"8851",
	145 => X"8296",
	146 => X"801A",
	147 => X"80EE",
	148 => X"850D",
	149 => X"8C5B",
	150 => X"96A8",
	151 => X"A3AF",
	152 => X"B31A",
	153 => X"C483",
	154 => X"D776",
	155 => X"EB76",
	156 => X"0000",
	157 => X"1488",
	158 => X"2888",
	159 => X"3B7B",
	160 => X"4CE4",
	161 => X"5C4F",
	162 => X"6956",
	163 => X"73A3",
	164 => X"7AF1",
	165 => X"7F10",
	166 => X"7FE4",
	167 => X"7D68",
	168 => X"77AD",
	169 => X"6ED9",
	170 => X"6325",
	171 => X"54E0",
	172 => X"4468",
	173 => X"322B",
	174 => X"1EA1",
	175 => X"0A4C",
	176 => X"F5B2",
	177 => X"E15D",
	178 => X"CDD3",
	179 => X"BB96",
	180 => X"AB1E",
	181 => X"9CD9",
	182 => X"9125",
	183 => X"8851",
	184 => X"8296",
	185 => X"801A",
	186 => X"80EE",
	187 => X"850D",
	188 => X"8C5B",
	189 => X"96A8",
	190 => X"A3AF",
	191 => X"B31A",
	192 => X"C483",
	193 => X"D776",
	194 => X"EB76",
	195 => X"0000",
	196 => X"1488",
	197 => X"2888",
	198 => X"3B7B",
	199 => X"4CE4",
	200 => X"5C4F",
	201 => X"6956",
	202 => X"73A3",
	203 => X"7AF1",
	204 => X"7F10",
	205 => X"7FE4",
	206 => X"7D68",
	207 => X"77AD",
	208 => X"6ED9",
	209 => X"6325",
	210 => X"54E0",
	211 => X"4468",
	212 => X"322B",
	213 => X"1EA1",
	214 => X"0A4C",
	215 => X"F5B2",
	216 => X"E15D",
	217 => X"CDD3",
	218 => X"BB96",
	219 => X"AB1E",
	220 => X"9CD9",
	221 => X"9125",
	222 => X"8851",
	223 => X"8296",
	224 => X"801A",
	225 => X"80EE",
	226 => X"850D",
	227 => X"8C5B",
	228 => X"96A8",
	229 => X"A3AF",
	230 => X"B31A",
	231 => X"C483",
	232 => X"D776",
	233 => X"EB76",
	234 => X"0000",
	235 => X"1488",
	236 => X"2888",
	237 => X"3B7B",
	238 => X"4CE4",
	239 => X"5C4F",
	240 => X"6956",
	241 => X"73A3",
	242 => X"7AF1",
	243 => X"7F10",
	244 => X"7FE4",
	245 => X"7D68",
	246 => X"77AD",
	247 => X"6ED9",
	others => X"0000"
);

CONSTANT A5: hex := (
	000 => X"0000",
	001 => X"15A1",
	002 => X"2AA3",
	003 => X"3E6C",
	004 => X"5068",
	005 => X"6015",
	006 => X"6CFE",
	007 => X"76C4",
	008 => X"7D1F",
	009 => X"7FE1",
	010 => X"7EF5",
	011 => X"7A62",
	012 => X"724A",
	013 => X"66E8",
	014 => X"5890",
	015 => X"47AC",
	016 => X"34B8",
	017 => X"2040",
	018 => X"0ADA",
	019 => X"F524",
	020 => X"DFBE",
	021 => X"CB46",
	022 => X"B852",
	023 => X"A76E",
	024 => X"9916",
	025 => X"8DB4",
	026 => X"859C",
	027 => X"8109",
	028 => X"801D",
	029 => X"82DF",
	030 => X"893A",
	031 => X"9300",
	032 => X"9FE9",
	033 => X"AF96",
	034 => X"C192",
	035 => X"D55B",
	036 => X"EA5D",
	037 => X"0000",
	038 => X"15A1",
	039 => X"2AA3",
	040 => X"3E6C",
	041 => X"5068",
	042 => X"6015",
	043 => X"6CFE",
	044 => X"76C4",
	045 => X"7D1F",
	046 => X"7FE1",
	047 => X"7EF5",
	048 => X"7A62",
	049 => X"724A",
	050 => X"66E8",
	051 => X"5890",
	052 => X"47AC",
	053 => X"34B8",
	054 => X"2040",
	055 => X"0ADA",
	056 => X"F524",
	057 => X"DFBE",
	058 => X"CB46",
	059 => X"B852",
	060 => X"A76E",
	061 => X"9916",
	062 => X"8DB4",
	063 => X"859C",
	064 => X"8109",
	065 => X"801D",
	066 => X"82DF",
	067 => X"893A",
	068 => X"9300",
	069 => X"9FE9",
	070 => X"AF96",
	071 => X"C192",
	072 => X"D55B",
	073 => X"EA5D",
	074 => X"FFFE",
	075 => X"15A1",
	076 => X"2AA3",
	077 => X"3E6C",
	078 => X"5068",
	079 => X"6015",
	080 => X"6CFE",
	081 => X"76C4",
	082 => X"7D1F",
	083 => X"7FE1",
	084 => X"7EF5",
	085 => X"7A62",
	086 => X"724A",
	087 => X"66E8",
	088 => X"5890",
	089 => X"47AC",
	090 => X"34B8",
	091 => X"2040",
	092 => X"0ADA",
	093 => X"F524",
	094 => X"DFBE",
	095 => X"CB46",
	096 => X"B852",
	097 => X"A76E",
	098 => X"9916",
	099 => X"8DB4",
	100 => X"859C",
	101 => X"8109",
	102 => X"801D",
	103 => X"82DF",
	104 => X"893A",
	105 => X"9300",
	106 => X"9FE9",
	107 => X"AF96",
	108 => X"C192",
	109 => X"D55B",
	110 => X"EA5D",
	111 => X"FFFE",
	112 => X"15A1",
	113 => X"2AA3",
	114 => X"3E6C",
	115 => X"5068",
	116 => X"6015",
	117 => X"6CFE",
	118 => X"76C4",
	119 => X"7D1F",
	120 => X"7FE1",
	121 => X"7EF5",
	122 => X"7A62",
	123 => X"724A",
	124 => X"66E8",
	125 => X"5890",
	126 => X"47AC",
	127 => X"34B8",
	128 => X"2040",
	129 => X"0ADA",
	130 => X"F524",
	131 => X"DFBE",
	132 => X"CB46",
	133 => X"B852",
	134 => X"A76E",
	135 => X"9916",
	136 => X"8DB4",
	137 => X"859C",
	138 => X"8109",
	139 => X"801D",
	140 => X"82DF",
	141 => X"893A",
	142 => X"9300",
	143 => X"9FE9",
	144 => X"AF96",
	145 => X"C192",
	146 => X"D55B",
	147 => X"EA5D",
	148 => X"0000",
	149 => X"15A1",
	150 => X"2AA3",
	151 => X"3E6C",
	152 => X"5068",
	153 => X"6015",
	154 => X"6CFE",
	155 => X"76C4",
	156 => X"7D1F",
	157 => X"7FE1",
	158 => X"7EF5",
	159 => X"7A62",
	160 => X"724A",
	161 => X"66E8",
	162 => X"5890",
	163 => X"47AC",
	164 => X"34B8",
	165 => X"2040",
	166 => X"0ADA",
	167 => X"F524",
	168 => X"DFBE",
	169 => X"CB46",
	170 => X"B852",
	171 => X"A76E",
	172 => X"9916",
	173 => X"8DB4",
	174 => X"859C",
	175 => X"8109",
	176 => X"801D",
	177 => X"82DF",
	178 => X"893A",
	179 => X"9300",
	180 => X"9FE9",
	181 => X"AF96",
	182 => X"C192",
	183 => X"D55B",
	184 => X"EA5D",
	185 => X"0000",
	186 => X"15A1",
	187 => X"2AA3",
	188 => X"3E6C",
	189 => X"5068",
	190 => X"6015",
	191 => X"6CFE",
	192 => X"76C4",
	193 => X"7D1F",
	194 => X"7FE1",
	195 => X"7EF5",
	196 => X"7A62",
	197 => X"724A",
	198 => X"66E8",
	199 => X"5890",
	200 => X"47AC",
	201 => X"34B8",
	202 => X"2040",
	203 => X"0ADA",
	204 => X"F524",
	205 => X"DFBE",
	206 => X"CB46",
	207 => X"B852",
	208 => X"A76E",
	209 => X"9916",
	210 => X"8DB4",
	211 => X"859C",
	212 => X"8109",
	213 => X"801D",
	214 => X"82DF",
	215 => X"893A",
	216 => X"9300",
	217 => X"9FE9",
	218 => X"AF96",
	219 => X"C192",
	220 => X"D55B",
	221 => X"EA5D",
	222 => X"0000",
	223 => X"15A1",
	224 => X"2AA3",
	225 => X"3E6C",
	226 => X"5068",
	227 => X"6015",
	228 => X"6CFE",
	229 => X"76C4",
	230 => X"7D1F",
	231 => X"7FE1",
	232 => X"7EF5",
	233 => X"7A62",
	234 => X"724A",
	235 => X"66E8",
	236 => X"5890",
	237 => X"47AC",
	238 => X"34B8",
	239 => X"2040",
	240 => X"0ADA",
	241 => X"F524",
	242 => X"DFBE",
	243 => X"CB46",
	244 => X"B852",
	245 => X"A76E",
	246 => X"9916",
	247 => X"8DB4",
	others => X"0000"
);

CONSTANT AS5: hex := (
	000 => X"0000",
	001 => X"16DA",
	002 => X"2CF9",
	003 => X"41A6",
	004 => X"5436",
	005 => X"6412",
	006 => X"70B6",
	007 => X"79BB",
	008 => X"7ED6",
	009 => X"7FDE",
	010 => X"7CC9",
	011 => X"75B2",
	012 => X"6AD2",
	013 => X"5C83",
	014 => X"4B3B",
	015 => X"3789",
	016 => X"220D",
	017 => X"0B79",
	018 => X"F485",
	019 => X"DDF1",
	020 => X"C875",
	021 => X"B4C3",
	022 => X"A37B",
	023 => X"952C",
	024 => X"8A4C",
	025 => X"8335",
	026 => X"8020",
	027 => X"8128",
	028 => X"8643",
	029 => X"8F48",
	030 => X"9BEC",
	031 => X"ABC8",
	032 => X"BE58",
	033 => X"D305",
	034 => X"E924",
	035 => X"FFFE",
	036 => X"16DA",
	037 => X"2CF9",
	038 => X"41A6",
	039 => X"5436",
	040 => X"6412",
	041 => X"70B6",
	042 => X"79BB",
	043 => X"7ED6",
	044 => X"7FDE",
	045 => X"7CC9",
	046 => X"75B2",
	047 => X"6AD2",
	048 => X"5C83",
	049 => X"4B3B",
	050 => X"3789",
	051 => X"220D",
	052 => X"0B79",
	053 => X"F485",
	054 => X"DDF1",
	055 => X"C875",
	056 => X"B4C3",
	057 => X"A37B",
	058 => X"952C",
	059 => X"8A4C",
	060 => X"8335",
	061 => X"8020",
	062 => X"8128",
	063 => X"8643",
	064 => X"8F48",
	065 => X"9BEC",
	066 => X"ABC8",
	067 => X"BE58",
	068 => X"D305",
	069 => X"E924",
	070 => X"0000",
	071 => X"16DA",
	072 => X"2CF9",
	073 => X"41A6",
	074 => X"5436",
	075 => X"6412",
	076 => X"70B6",
	077 => X"79BB",
	078 => X"7ED6",
	079 => X"7FDE",
	080 => X"7CC9",
	081 => X"75B2",
	082 => X"6AD2",
	083 => X"5C83",
	084 => X"4B3B",
	085 => X"3789",
	086 => X"220D",
	087 => X"0B79",
	088 => X"F485",
	089 => X"DDF1",
	090 => X"C875",
	091 => X"B4C3",
	092 => X"A37B",
	093 => X"952C",
	094 => X"8A4C",
	095 => X"8335",
	096 => X"8020",
	097 => X"8128",
	098 => X"8643",
	099 => X"8F48",
	100 => X"9BEC",
	101 => X"ABC8",
	102 => X"BE58",
	103 => X"D305",
	104 => X"E924",
	105 => X"0000",
	106 => X"16DA",
	107 => X"2CF9",
	108 => X"41A6",
	109 => X"5436",
	110 => X"6412",
	111 => X"70B6",
	112 => X"79BB",
	113 => X"7ED6",
	114 => X"7FDE",
	115 => X"7CC9",
	116 => X"75B2",
	117 => X"6AD2",
	118 => X"5C83",
	119 => X"4B3B",
	120 => X"3789",
	121 => X"220D",
	122 => X"0B79",
	123 => X"F485",
	124 => X"DDF1",
	125 => X"C875",
	126 => X"B4C3",
	127 => X"A37B",
	128 => X"952C",
	129 => X"8A4C",
	130 => X"8335",
	131 => X"8020",
	132 => X"8128",
	133 => X"8643",
	134 => X"8F48",
	135 => X"9BEC",
	136 => X"ABC8",
	137 => X"BE58",
	138 => X"D305",
	139 => X"E924",
	140 => X"FFFE",
	141 => X"16DA",
	142 => X"2CF9",
	143 => X"41A6",
	144 => X"5436",
	145 => X"6412",
	146 => X"70B6",
	147 => X"79BB",
	148 => X"7ED6",
	149 => X"7FDE",
	150 => X"7CC9",
	151 => X"75B2",
	152 => X"6AD2",
	153 => X"5C83",
	154 => X"4B3B",
	155 => X"3789",
	156 => X"220D",
	157 => X"0B79",
	158 => X"F485",
	159 => X"DDF1",
	160 => X"C875",
	161 => X"B4C3",
	162 => X"A37B",
	163 => X"952C",
	164 => X"8A4C",
	165 => X"8335",
	166 => X"8020",
	167 => X"8128",
	168 => X"8643",
	169 => X"8F48",
	170 => X"9BEC",
	171 => X"ABC8",
	172 => X"BE58",
	173 => X"D305",
	174 => X"E924",
	175 => X"FFFE",
	176 => X"16DA",
	177 => X"2CF9",
	178 => X"41A6",
	179 => X"5436",
	180 => X"6412",
	181 => X"70B6",
	182 => X"79BB",
	183 => X"7ED6",
	184 => X"7FDE",
	185 => X"7CC9",
	186 => X"75B2",
	187 => X"6AD2",
	188 => X"5C83",
	189 => X"4B3B",
	190 => X"3789",
	191 => X"220D",
	192 => X"0B79",
	193 => X"F485",
	194 => X"DDF1",
	195 => X"C875",
	196 => X"B4C3",
	197 => X"A37B",
	198 => X"952C",
	199 => X"8A4C",
	200 => X"8335",
	201 => X"8020",
	202 => X"8128",
	203 => X"8643",
	204 => X"8F48",
	205 => X"9BEC",
	206 => X"ABC8",
	207 => X"BE58",
	208 => X"D305",
	209 => X"E924",
	210 => X"FFFE",
	211 => X"16DA",
	212 => X"2CF9",
	213 => X"41A6",
	214 => X"5436",
	215 => X"6412",
	216 => X"70B6",
	217 => X"79BB",
	218 => X"7ED6",
	219 => X"7FDE",
	220 => X"7CC9",
	221 => X"75B2",
	222 => X"6AD2",
	223 => X"5C83",
	224 => X"4B3B",
	225 => X"3789",
	226 => X"220D",
	227 => X"0B79",
	228 => X"F485",
	229 => X"DDF1",
	230 => X"C875",
	231 => X"B4C3",
	232 => X"A37B",
	233 => X"952C",
	234 => X"8A4C",
	235 => X"8335",
	236 => X"8020",
	237 => X"8128",
	238 => X"8643",
	239 => X"8F48",
	240 => X"9BEC",
	241 => X"ABC8",
	242 => X"BE58",
	243 => X"D305",
	244 => X"E924",
	245 => X"FFFE",
	246 => X"16DA",
	247 => X"2CF9",
	others => X"0000"
);

CONSTANT B5: hex := (
	000 => X"0000",
	001 => X"1839",
	002 => X"2F92",
	003 => X"4533",
	004 => X"5853",
	005 => X"6843",
	006 => X"746D",
	007 => X"7C63",
	008 => X"7FD9",
	009 => X"7EB1",
	010 => X"78F4",
	011 => X"6ED9",
	012 => X"60BB",
	013 => X"4F1F",
	014 => X"3AA6",
	015 => X"240F",
	016 => X"0C2A",
	017 => X"F3D4",
	018 => X"DBEF",
	019 => X"C558",
	020 => X"B0DF",
	021 => X"9F43",
	022 => X"9125",
	023 => X"870A",
	024 => X"814D",
	025 => X"8025",
	026 => X"839B",
	027 => X"8B91",
	028 => X"97BB",
	029 => X"A7AB",
	030 => X"BACB",
	031 => X"D06C",
	032 => X"E7C5",
	033 => X"0000",
	034 => X"1839",
	035 => X"2F92",
	036 => X"4533",
	037 => X"5853",
	038 => X"6843",
	039 => X"746D",
	040 => X"7C63",
	041 => X"7FD9",
	042 => X"7EB1",
	043 => X"78F4",
	044 => X"6ED9",
	045 => X"60BB",
	046 => X"4F1F",
	047 => X"3AA6",
	048 => X"240F",
	049 => X"0C2A",
	050 => X"F3D4",
	051 => X"DBEF",
	052 => X"C558",
	053 => X"B0DF",
	054 => X"9F43",
	055 => X"9125",
	056 => X"870A",
	057 => X"814D",
	058 => X"8025",
	059 => X"839B",
	060 => X"8B91",
	061 => X"97BB",
	062 => X"A7AB",
	063 => X"BACB",
	064 => X"D06C",
	065 => X"E7C5",
	066 => X"FFFE",
	067 => X"1839",
	068 => X"2F92",
	069 => X"4533",
	070 => X"5853",
	071 => X"6843",
	072 => X"746D",
	073 => X"7C63",
	074 => X"7FD9",
	075 => X"7EB1",
	076 => X"78F4",
	077 => X"6ED9",
	078 => X"60BB",
	079 => X"4F1F",
	080 => X"3AA6",
	081 => X"240F",
	082 => X"0C2A",
	083 => X"F3D4",
	084 => X"DBEF",
	085 => X"C558",
	086 => X"B0DF",
	087 => X"9F43",
	088 => X"9125",
	089 => X"870A",
	090 => X"814D",
	091 => X"8025",
	092 => X"839B",
	093 => X"8B91",
	094 => X"97BB",
	095 => X"A7AB",
	096 => X"BACB",
	097 => X"D06C",
	098 => X"E7C5",
	099 => X"FFFE",
	100 => X"1839",
	101 => X"2F92",
	102 => X"4533",
	103 => X"5853",
	104 => X"6843",
	105 => X"746D",
	106 => X"7C63",
	107 => X"7FD9",
	108 => X"7EB1",
	109 => X"78F4",
	110 => X"6ED9",
	111 => X"60BB",
	112 => X"4F1F",
	113 => X"3AA6",
	114 => X"240F",
	115 => X"0C2A",
	116 => X"F3D4",
	117 => X"DBEF",
	118 => X"C558",
	119 => X"B0DF",
	120 => X"9F43",
	121 => X"9125",
	122 => X"870A",
	123 => X"814D",
	124 => X"8025",
	125 => X"839B",
	126 => X"8B91",
	127 => X"97BB",
	128 => X"A7AB",
	129 => X"BACB",
	130 => X"D06C",
	131 => X"E7C5",
	132 => X"0000",
	133 => X"1839",
	134 => X"2F92",
	135 => X"4533",
	136 => X"5853",
	137 => X"6843",
	138 => X"746D",
	139 => X"7C63",
	140 => X"7FD9",
	141 => X"7EB1",
	142 => X"78F4",
	143 => X"6ED9",
	144 => X"60BB",
	145 => X"4F1F",
	146 => X"3AA6",
	147 => X"240F",
	148 => X"0C2A",
	149 => X"F3D4",
	150 => X"DBEF",
	151 => X"C558",
	152 => X"B0DF",
	153 => X"9F43",
	154 => X"9125",
	155 => X"870A",
	156 => X"814D",
	157 => X"8025",
	158 => X"839B",
	159 => X"8B91",
	160 => X"97BB",
	161 => X"A7AB",
	162 => X"BACB",
	163 => X"D06C",
	164 => X"E7C5",
	165 => X"0000",
	166 => X"1839",
	167 => X"2F92",
	168 => X"4533",
	169 => X"5853",
	170 => X"6843",
	171 => X"746D",
	172 => X"7C63",
	173 => X"7FD9",
	174 => X"7EB1",
	175 => X"78F4",
	176 => X"6ED9",
	177 => X"60BB",
	178 => X"4F1F",
	179 => X"3AA6",
	180 => X"240F",
	181 => X"0C2A",
	182 => X"F3D4",
	183 => X"DBEF",
	184 => X"C558",
	185 => X"B0DF",
	186 => X"9F43",
	187 => X"9125",
	188 => X"870A",
	189 => X"814D",
	190 => X"8025",
	191 => X"839B",
	192 => X"8B91",
	193 => X"97BB",
	194 => X"A7AB",
	195 => X"BACB",
	196 => X"D06C",
	197 => X"E7C5",
	198 => X"0000",
	199 => X"1839",
	200 => X"2F92",
	201 => X"4533",
	202 => X"5853",
	203 => X"6843",
	204 => X"746D",
	205 => X"7C63",
	206 => X"7FD9",
	207 => X"7EB1",
	208 => X"78F4",
	209 => X"6ED9",
	210 => X"60BB",
	211 => X"4F1F",
	212 => X"3AA6",
	213 => X"240F",
	214 => X"0C2A",
	215 => X"F3D4",
	216 => X"DBEF",
	217 => X"C558",
	218 => X"B0DF",
	219 => X"9F43",
	220 => X"9125",
	221 => X"870A",
	222 => X"814D",
	223 => X"8025",
	224 => X"839B",
	225 => X"8B91",
	226 => X"97BB",
	227 => X"A7AB",
	228 => X"BACB",
	229 => X"D06C",
	230 => X"E7C5",
	231 => X"0000",
	232 => X"1839",
	233 => X"2F92",
	234 => X"4533",
	235 => X"5853",
	236 => X"6843",
	237 => X"746D",
	238 => X"7C63",
	239 => X"7FD9",
	240 => X"7EB1",
	241 => X"78F4",
	242 => X"6ED9",
	243 => X"60BB",
	244 => X"4F1F",
	245 => X"3AA6",
	246 => X"240F",
	247 => X"0C2A",
	others => X"0000"
);

CONSTANT C6: hex := (
	000 => X"0000",
	001 => X"19C3",
	002 => X"3279",
	003 => X"491E",
	004 => X"5CC5",
	005 => X"6C9F",
	006 => X"7807",
	007 => X"7E85",
	008 => X"7FD4",
	009 => X"7BE8",
	010 => X"72EA",
	011 => X"6537",
	012 => X"535F",
	013 => X"3E1D",
	014 => X"2651",
	015 => X"0CF2",
	016 => X"F30C",
	017 => X"D9AD",
	018 => X"C1E1",
	019 => X"AC9F",
	020 => X"9AC7",
	021 => X"8D14",
	022 => X"8416",
	023 => X"802A",
	024 => X"8179",
	025 => X"87F7",
	026 => X"935F",
	027 => X"A339",
	028 => X"B6E0",
	029 => X"CD85",
	030 => X"E63B",
	031 => X"0000",
	032 => X"19C3",
	033 => X"3279",
	034 => X"491E",
	035 => X"5CC5",
	036 => X"6C9F",
	037 => X"7807",
	038 => X"7E85",
	039 => X"7FD4",
	040 => X"7BE8",
	041 => X"72EA",
	042 => X"6537",
	043 => X"535F",
	044 => X"3E1D",
	045 => X"2651",
	046 => X"0CF2",
	047 => X"F30C",
	048 => X"D9AD",
	049 => X"C1E1",
	050 => X"AC9F",
	051 => X"9AC7",
	052 => X"8D14",
	053 => X"8416",
	054 => X"802A",
	055 => X"8179",
	056 => X"87F7",
	057 => X"935F",
	058 => X"A339",
	059 => X"B6E0",
	060 => X"CD85",
	061 => X"E63B",
	062 => X"0000",
	063 => X"19C3",
	064 => X"3279",
	065 => X"491E",
	066 => X"5CC5",
	067 => X"6C9F",
	068 => X"7807",
	069 => X"7E85",
	070 => X"7FD4",
	071 => X"7BE8",
	072 => X"72EA",
	073 => X"6537",
	074 => X"535F",
	075 => X"3E1D",
	076 => X"2651",
	077 => X"0CF2",
	078 => X"F30C",
	079 => X"D9AD",
	080 => X"C1E1",
	081 => X"AC9F",
	082 => X"9AC7",
	083 => X"8D14",
	084 => X"8416",
	085 => X"802A",
	086 => X"8179",
	087 => X"87F7",
	088 => X"935F",
	089 => X"A339",
	090 => X"B6E0",
	091 => X"CD85",
	092 => X"E63B",
	093 => X"0000",
	094 => X"19C3",
	095 => X"3279",
	096 => X"491E",
	097 => X"5CC5",
	098 => X"6C9F",
	099 => X"7807",
	100 => X"7E85",
	101 => X"7FD4",
	102 => X"7BE8",
	103 => X"72EA",
	104 => X"6537",
	105 => X"535F",
	106 => X"3E1D",
	107 => X"2651",
	108 => X"0CF2",
	109 => X"F30C",
	110 => X"D9AD",
	111 => X"C1E1",
	112 => X"AC9F",
	113 => X"9AC7",
	114 => X"8D14",
	115 => X"8416",
	116 => X"802A",
	117 => X"8179",
	118 => X"87F7",
	119 => X"935F",
	120 => X"A339",
	121 => X"B6E0",
	122 => X"CD85",
	123 => X"E63B",
	124 => X"FFFE",
	125 => X"19C3",
	126 => X"3279",
	127 => X"491E",
	128 => X"5CC5",
	129 => X"6C9F",
	130 => X"7807",
	131 => X"7E85",
	132 => X"7FD4",
	133 => X"7BE8",
	134 => X"72EA",
	135 => X"6537",
	136 => X"535F",
	137 => X"3E1D",
	138 => X"2651",
	139 => X"0CF2",
	140 => X"F30C",
	141 => X"D9AD",
	142 => X"C1E1",
	143 => X"AC9F",
	144 => X"9AC7",
	145 => X"8D14",
	146 => X"8416",
	147 => X"802A",
	148 => X"8179",
	149 => X"87F7",
	150 => X"935F",
	151 => X"A339",
	152 => X"B6E0",
	153 => X"CD85",
	154 => X"E63B",
	155 => X"FFFE",
	156 => X"19C3",
	157 => X"3279",
	158 => X"491E",
	159 => X"5CC5",
	160 => X"6C9F",
	161 => X"7807",
	162 => X"7E85",
	163 => X"7FD4",
	164 => X"7BE8",
	165 => X"72EA",
	166 => X"6537",
	167 => X"535F",
	168 => X"3E1D",
	169 => X"2651",
	170 => X"0CF2",
	171 => X"F30C",
	172 => X"D9AD",
	173 => X"C1E1",
	174 => X"AC9F",
	175 => X"9AC7",
	176 => X"8D14",
	177 => X"8416",
	178 => X"802A",
	179 => X"8179",
	180 => X"87F7",
	181 => X"935F",
	182 => X"A339",
	183 => X"B6E0",
	184 => X"CD85",
	185 => X"E63B",
	186 => X"FFFE",
	187 => X"19C3",
	188 => X"3279",
	189 => X"491E",
	190 => X"5CC5",
	191 => X"6C9F",
	192 => X"7807",
	193 => X"7E85",
	194 => X"7FD4",
	195 => X"7BE8",
	196 => X"72EA",
	197 => X"6537",
	198 => X"535F",
	199 => X"3E1D",
	200 => X"2651",
	201 => X"0CF2",
	202 => X"F30C",
	203 => X"D9AD",
	204 => X"C1E1",
	205 => X"AC9F",
	206 => X"9AC7",
	207 => X"8D14",
	208 => X"8416",
	209 => X"802A",
	210 => X"8179",
	211 => X"87F7",
	212 => X"935F",
	213 => X"A339",
	214 => X"B6E0",
	215 => X"CD85",
	216 => X"E63B",
	217 => X"FFFE",
	218 => X"19C3",
	219 => X"3279",
	220 => X"491E",
	221 => X"5CC5",
	222 => X"6C9F",
	223 => X"7807",
	224 => X"7E85",
	225 => X"7FD4",
	226 => X"7BE8",
	227 => X"72EA",
	228 => X"6537",
	229 => X"535F",
	230 => X"3E1D",
	231 => X"2651",
	232 => X"0CF2",
	233 => X"F30C",
	234 => X"D9AD",
	235 => X"C1E1",
	236 => X"AC9F",
	237 => X"9AC7",
	238 => X"8D14",
	239 => X"8416",
	240 => X"802A",
	241 => X"8179",
	242 => X"87F7",
	243 => X"935F",
	244 => X"A339",
	245 => X"B6E0",
	246 => X"CD85",
	247 => X"E63B",
	others => X"0000"
);

CONSTANT CS6: hex := (
	000 => X"0000",
	001 => X"1B83",
	002 => X"35BE",
	003 => X"4D75",
	004 => X"618D",
	005 => X"7116",
	006 => X"7B54",
	007 => X"7FCE",
	008 => X"7E4F",
	009 => X"76E7",
	010 => X"69F0",
	011 => X"5805",
	012 => X"41FD",
	013 => X"28DE",
	014 => X"0DD6",
	015 => X"F228",
	016 => X"D720",
	017 => X"BE01",
	018 => X"A7F9",
	019 => X"960E",
	020 => X"8917",
	021 => X"81AF",
	022 => X"8030",
	023 => X"84AA",
	024 => X"8EE8",
	025 => X"9E71",
	026 => X"B289",
	027 => X"CA40",
	028 => X"E47B",
	029 => X"FFFE",
	030 => X"1B83",
	031 => X"35BE",
	032 => X"4D75",
	033 => X"618D",
	034 => X"7116",
	035 => X"7B54",
	036 => X"7FCE",
	037 => X"7E4F",
	038 => X"76E7",
	039 => X"69F0",
	040 => X"5805",
	041 => X"41FD",
	042 => X"28DE",
	043 => X"0DD6",
	044 => X"F228",
	045 => X"D720",
	046 => X"BE01",
	047 => X"A7F9",
	048 => X"960E",
	049 => X"8917",
	050 => X"81AF",
	051 => X"8030",
	052 => X"84AA",
	053 => X"8EE8",
	054 => X"9E71",
	055 => X"B289",
	056 => X"CA40",
	057 => X"E47B",
	058 => X"FFFE",
	059 => X"1B83",
	060 => X"35BE",
	061 => X"4D75",
	062 => X"618D",
	063 => X"7116",
	064 => X"7B54",
	065 => X"7FCE",
	066 => X"7E4F",
	067 => X"76E7",
	068 => X"69F0",
	069 => X"5805",
	070 => X"41FD",
	071 => X"28DE",
	072 => X"0DD6",
	073 => X"F228",
	074 => X"D720",
	075 => X"BE01",
	076 => X"A7F9",
	077 => X"960E",
	078 => X"8917",
	079 => X"81AF",
	080 => X"8030",
	081 => X"84AA",
	082 => X"8EE8",
	083 => X"9E71",
	084 => X"B289",
	085 => X"CA40",
	086 => X"E47B",
	087 => X"FFFE",
	088 => X"1B83",
	089 => X"35BE",
	090 => X"4D75",
	091 => X"618D",
	092 => X"7116",
	093 => X"7B54",
	094 => X"7FCE",
	095 => X"7E4F",
	096 => X"76E7",
	097 => X"69F0",
	098 => X"5805",
	099 => X"41FD",
	100 => X"28DE",
	101 => X"0DD6",
	102 => X"F228",
	103 => X"D720",
	104 => X"BE01",
	105 => X"A7F9",
	106 => X"960E",
	107 => X"8917",
	108 => X"81AF",
	109 => X"8030",
	110 => X"84AA",
	111 => X"8EE8",
	112 => X"9E71",
	113 => X"B289",
	114 => X"CA40",
	115 => X"E47B",
	116 => X"0000",
	117 => X"1B83",
	118 => X"35BE",
	119 => X"4D75",
	120 => X"618D",
	121 => X"7116",
	122 => X"7B54",
	123 => X"7FCE",
	124 => X"7E4F",
	125 => X"76E7",
	126 => X"69F0",
	127 => X"5805",
	128 => X"41FD",
	129 => X"28DE",
	130 => X"0DD6",
	131 => X"F228",
	132 => X"D720",
	133 => X"BE01",
	134 => X"A7F9",
	135 => X"960E",
	136 => X"8917",
	137 => X"81AF",
	138 => X"8030",
	139 => X"84AA",
	140 => X"8EE8",
	141 => X"9E71",
	142 => X"B289",
	143 => X"CA40",
	144 => X"E47B",
	145 => X"0000",
	146 => X"1B83",
	147 => X"35BE",
	148 => X"4D75",
	149 => X"618D",
	150 => X"7116",
	151 => X"7B54",
	152 => X"7FCE",
	153 => X"7E4F",
	154 => X"76E7",
	155 => X"69F0",
	156 => X"5805",
	157 => X"41FD",
	158 => X"28DE",
	159 => X"0DD6",
	160 => X"F228",
	161 => X"D720",
	162 => X"BE01",
	163 => X"A7F9",
	164 => X"960E",
	165 => X"8917",
	166 => X"81AF",
	167 => X"8030",
	168 => X"84AA",
	169 => X"8EE8",
	170 => X"9E71",
	171 => X"B289",
	172 => X"CA40",
	173 => X"E47B",
	174 => X"0000",
	175 => X"1B83",
	176 => X"35BE",
	177 => X"4D75",
	178 => X"618D",
	179 => X"7116",
	180 => X"7B54",
	181 => X"7FCE",
	182 => X"7E4F",
	183 => X"76E7",
	184 => X"69F0",
	185 => X"5805",
	186 => X"41FD",
	187 => X"28DE",
	188 => X"0DD6",
	189 => X"F228",
	190 => X"D720",
	191 => X"BE01",
	192 => X"A7F9",
	193 => X"960E",
	194 => X"8917",
	195 => X"81AF",
	196 => X"8030",
	197 => X"84AA",
	198 => X"8EE8",
	199 => X"9E71",
	200 => X"B289",
	201 => X"CA40",
	202 => X"E47B",
	203 => X"0000",
	204 => X"1B83",
	205 => X"35BE",
	206 => X"4D75",
	207 => X"618D",
	208 => X"7116",
	209 => X"7B54",
	210 => X"7FCE",
	211 => X"7E4F",
	212 => X"76E7",
	213 => X"69F0",
	214 => X"5805",
	215 => X"41FD",
	216 => X"28DE",
	217 => X"0DD6",
	218 => X"F228",
	219 => X"D720",
	220 => X"BE01",
	221 => X"A7F9",
	222 => X"960E",
	223 => X"8917",
	224 => X"81AF",
	225 => X"8030",
	226 => X"84AA",
	227 => X"8EE8",
	228 => X"9E71",
	229 => X"B289",
	230 => X"CA40",
	231 => X"E47B",
	232 => X"0000",
	233 => X"1B83",
	234 => X"35BE",
	235 => X"4D75",
	236 => X"618D",
	237 => X"7116",
	238 => X"7B54",
	239 => X"7FCE",
	240 => X"7E4F",
	241 => X"76E7",
	242 => X"69F0",
	243 => X"5805",
	244 => X"41FD",
	245 => X"28DE",
	246 => X"0DD6",
	247 => X"F228",
	others => X"0000"
);

CONSTANT D6: hex := (
	000 => X"0000",
	001 => X"1C7B",
	002 => X"3789",
	003 => X"4FCD",
	004 => X"6412",
	005 => X"7352",
	006 => X"7CC9",
	007 => X"7FFF",
	008 => X"7CC9",
	009 => X"7352",
	010 => X"6412",
	011 => X"4FCD",
	012 => X"3789",
	013 => X"1C7B",
	014 => X"FFFE",
	015 => X"E383",
	016 => X"C875",
	017 => X"B031",
	018 => X"9BEC",
	019 => X"8CAC",
	020 => X"8335",
	021 => X"8000",
	022 => X"8335",
	023 => X"8CAC",
	024 => X"9BEC",
	025 => X"B031",
	026 => X"C875",
	027 => X"E383",
	028 => X"FFFE",
	029 => X"1C7B",
	030 => X"3789",
	031 => X"4FCD",
	032 => X"6412",
	033 => X"7352",
	034 => X"7CC9",
	035 => X"7FFF",
	036 => X"7CC9",
	037 => X"7352",
	038 => X"6412",
	039 => X"4FCD",
	040 => X"3789",
	041 => X"1C7B",
	042 => X"0000",
	043 => X"E383",
	044 => X"C875",
	045 => X"B031",
	046 => X"9BEC",
	047 => X"8CAC",
	048 => X"8335",
	049 => X"8000",
	050 => X"8335",
	051 => X"8CAC",
	052 => X"9BEC",
	053 => X"B031",
	054 => X"C875",
	055 => X"E383",
	056 => X"0000",
	057 => X"1C7B",
	058 => X"3789",
	059 => X"4FCD",
	060 => X"6412",
	061 => X"7352",
	062 => X"7CC9",
	063 => X"7FFF",
	064 => X"7CC9",
	065 => X"7352",
	066 => X"6412",
	067 => X"4FCD",
	068 => X"3789",
	069 => X"1C7B",
	070 => X"FFFE",
	071 => X"E383",
	072 => X"C875",
	073 => X"B031",
	074 => X"9BEC",
	075 => X"8CAC",
	076 => X"8335",
	077 => X"8000",
	078 => X"8335",
	079 => X"8CAC",
	080 => X"9BEC",
	081 => X"B031",
	082 => X"C875",
	083 => X"E383",
	084 => X"0000",
	085 => X"1C7B",
	086 => X"3789",
	087 => X"4FCD",
	088 => X"6412",
	089 => X"7352",
	090 => X"7CC9",
	091 => X"7FFF",
	092 => X"7CC9",
	093 => X"7352",
	094 => X"6412",
	095 => X"4FCD",
	096 => X"3789",
	097 => X"1C7B",
	098 => X"FFFE",
	099 => X"E383",
	100 => X"C875",
	101 => X"B031",
	102 => X"9BEC",
	103 => X"8CAC",
	104 => X"8335",
	105 => X"8000",
	106 => X"8335",
	107 => X"8CAC",
	108 => X"9BEC",
	109 => X"B031",
	110 => X"C875",
	111 => X"E383",
	112 => X"0000",
	113 => X"1C7B",
	114 => X"3789",
	115 => X"4FCD",
	116 => X"6412",
	117 => X"7352",
	118 => X"7CC9",
	119 => X"7FFF",
	120 => X"7CC9",
	121 => X"7352",
	122 => X"6412",
	123 => X"4FCD",
	124 => X"3789",
	125 => X"1C7B",
	126 => X"FFFE",
	127 => X"E383",
	128 => X"C875",
	129 => X"B031",
	130 => X"9BEC",
	131 => X"8CAC",
	132 => X"8335",
	133 => X"8000",
	134 => X"8335",
	135 => X"8CAC",
	136 => X"9BEC",
	137 => X"B031",
	138 => X"C875",
	139 => X"E383",
	140 => X"0000",
	141 => X"1C7B",
	142 => X"3789",
	143 => X"4FCD",
	144 => X"6412",
	145 => X"7352",
	146 => X"7CC9",
	147 => X"7FFF",
	148 => X"7CC9",
	149 => X"7352",
	150 => X"6412",
	151 => X"4FCD",
	152 => X"3789",
	153 => X"1C7B",
	154 => X"FFFE",
	155 => X"E383",
	156 => X"C875",
	157 => X"B031",
	158 => X"9BEC",
	159 => X"8CAC",
	160 => X"8335",
	161 => X"8000",
	162 => X"8335",
	163 => X"8CAC",
	164 => X"9BEC",
	165 => X"B031",
	166 => X"C875",
	167 => X"E383",
	168 => X"0000",
	169 => X"1C7B",
	170 => X"3789",
	171 => X"4FCD",
	172 => X"6412",
	173 => X"7352",
	174 => X"7CC9",
	175 => X"7FFF",
	176 => X"7CC9",
	177 => X"7352",
	178 => X"6412",
	179 => X"4FCD",
	180 => X"3789",
	181 => X"1C7B",
	182 => X"0000",
	183 => X"E383",
	184 => X"C875",
	185 => X"B031",
	186 => X"9BEC",
	187 => X"8CAC",
	188 => X"8335",
	189 => X"8000",
	190 => X"8335",
	191 => X"8CAC",
	192 => X"9BEC",
	193 => X"B031",
	194 => X"C875",
	195 => X"E383",
	196 => X"FFFE",
	197 => X"1C7B",
	198 => X"3789",
	199 => X"4FCD",
	200 => X"6412",
	201 => X"7352",
	202 => X"7CC9",
	203 => X"7FFF",
	204 => X"7CC9",
	205 => X"7352",
	206 => X"6412",
	207 => X"4FCD",
	208 => X"3789",
	209 => X"1C7B",
	210 => X"0000",
	211 => X"E383",
	212 => X"C875",
	213 => X"B031",
	214 => X"9BEC",
	215 => X"8CAC",
	216 => X"8335",
	217 => X"8000",
	218 => X"8335",
	219 => X"8CAC",
	220 => X"9BEC",
	221 => X"B031",
	222 => X"C875",
	223 => X"E383",
	224 => X"FFFE",
	225 => X"1C7B",
	226 => X"3789",
	227 => X"4FCD",
	228 => X"6412",
	229 => X"7352",
	230 => X"7CC9",
	231 => X"7FFF",
	232 => X"7CC9",
	233 => X"7352",
	234 => X"6412",
	235 => X"4FCD",
	236 => X"3789",
	237 => X"1C7B",
	238 => X"0000",
	239 => X"E383",
	240 => X"C875",
	241 => X"B031",
	242 => X"9BEC",
	243 => X"8CAC",
	244 => X"8335",
	245 => X"8000",
	246 => X"8335",
	247 => X"8CAC",
	others => X"0000"
);

CONSTANT DS6: hex := (
	000 => X"0000",
	001 => X"1EA1",
	002 => X"3B7B",
	003 => X"54E0",
	004 => X"6956",
	005 => X"77AD",
	006 => X"7F10",
	007 => X"7F10",
	008 => X"77AD",
	009 => X"6956",
	010 => X"54E0",
	011 => X"3B7B",
	012 => X"1EA1",
	013 => X"0000",
	014 => X"E15D",
	015 => X"C483",
	016 => X"AB1E",
	017 => X"96A8",
	018 => X"8851",
	019 => X"80EE",
	020 => X"80EE",
	021 => X"8851",
	022 => X"96A8",
	023 => X"AB1E",
	024 => X"C483",
	025 => X"E15D",
	026 => X"0000",
	027 => X"1EA1",
	028 => X"3B7B",
	029 => X"54E0",
	030 => X"6956",
	031 => X"77AD",
	032 => X"7F10",
	033 => X"7F10",
	034 => X"77AD",
	035 => X"6956",
	036 => X"54E0",
	037 => X"3B7B",
	038 => X"1EA1",
	039 => X"FFFE",
	040 => X"E15D",
	041 => X"C483",
	042 => X"AB1E",
	043 => X"96A8",
	044 => X"8851",
	045 => X"80EE",
	046 => X"80EE",
	047 => X"8851",
	048 => X"96A8",
	049 => X"AB1E",
	050 => X"C483",
	051 => X"E15D",
	052 => X"FFFE",
	053 => X"1EA1",
	054 => X"3B7B",
	055 => X"54E0",
	056 => X"6956",
	057 => X"77AD",
	058 => X"7F10",
	059 => X"7F10",
	060 => X"77AD",
	061 => X"6956",
	062 => X"54E0",
	063 => X"3B7B",
	064 => X"1EA1",
	065 => X"0000",
	066 => X"E15D",
	067 => X"C483",
	068 => X"AB1E",
	069 => X"96A8",
	070 => X"8851",
	071 => X"80EE",
	072 => X"80EE",
	073 => X"8851",
	074 => X"96A8",
	075 => X"AB1E",
	076 => X"C483",
	077 => X"E15D",
	078 => X"FFFE",
	079 => X"1EA1",
	080 => X"3B7B",
	081 => X"54E0",
	082 => X"6956",
	083 => X"77AD",
	084 => X"7F10",
	085 => X"7F10",
	086 => X"77AD",
	087 => X"6956",
	088 => X"54E0",
	089 => X"3B7B",
	090 => X"1EA1",
	091 => X"0000",
	092 => X"E15D",
	093 => X"C483",
	094 => X"AB1E",
	095 => X"96A8",
	096 => X"8851",
	097 => X"80EE",
	098 => X"80EE",
	099 => X"8851",
	100 => X"96A8",
	101 => X"AB1E",
	102 => X"C483",
	103 => X"E15D",
	104 => X"FFFE",
	105 => X"1EA1",
	106 => X"3B7B",
	107 => X"54E0",
	108 => X"6956",
	109 => X"77AD",
	110 => X"7F10",
	111 => X"7F10",
	112 => X"77AD",
	113 => X"6956",
	114 => X"54E0",
	115 => X"3B7B",
	116 => X"1EA1",
	117 => X"0000",
	118 => X"E15D",
	119 => X"C483",
	120 => X"AB1E",
	121 => X"96A8",
	122 => X"8851",
	123 => X"80EE",
	124 => X"80EE",
	125 => X"8851",
	126 => X"96A8",
	127 => X"AB1E",
	128 => X"C483",
	129 => X"E15D",
	130 => X"FFFE",
	131 => X"1EA1",
	132 => X"3B7B",
	133 => X"54E0",
	134 => X"6956",
	135 => X"77AD",
	136 => X"7F10",
	137 => X"7F10",
	138 => X"77AD",
	139 => X"6956",
	140 => X"54E0",
	141 => X"3B7B",
	142 => X"1EA1",
	143 => X"0000",
	144 => X"E15D",
	145 => X"C483",
	146 => X"AB1E",
	147 => X"96A8",
	148 => X"8851",
	149 => X"80EE",
	150 => X"80EE",
	151 => X"8851",
	152 => X"96A8",
	153 => X"AB1E",
	154 => X"C483",
	155 => X"E15D",
	156 => X"FFFE",
	157 => X"1EA1",
	158 => X"3B7B",
	159 => X"54E0",
	160 => X"6956",
	161 => X"77AD",
	162 => X"7F10",
	163 => X"7F10",
	164 => X"77AD",
	165 => X"6956",
	166 => X"54E0",
	167 => X"3B7B",
	168 => X"1EA1",
	169 => X"0000",
	170 => X"E15D",
	171 => X"C483",
	172 => X"AB1E",
	173 => X"96A8",
	174 => X"8851",
	175 => X"80EE",
	176 => X"80EE",
	177 => X"8851",
	178 => X"96A8",
	179 => X"AB1E",
	180 => X"C483",
	181 => X"E15D",
	182 => X"FFFE",
	183 => X"1EA1",
	184 => X"3B7B",
	185 => X"54E0",
	186 => X"6956",
	187 => X"77AD",
	188 => X"7F10",
	189 => X"7F10",
	190 => X"77AD",
	191 => X"6956",
	192 => X"54E0",
	193 => X"3B7B",
	194 => X"1EA1",
	195 => X"0000",
	196 => X"E15D",
	197 => X"C483",
	198 => X"AB1E",
	199 => X"96A8",
	200 => X"8851",
	201 => X"80EE",
	202 => X"80EE",
	203 => X"8851",
	204 => X"96A8",
	205 => X"AB1E",
	206 => X"C483",
	207 => X"E15D",
	208 => X"FFFE",
	209 => X"1EA1",
	210 => X"3B7B",
	211 => X"54E0",
	212 => X"6956",
	213 => X"77AD",
	214 => X"7F10",
	215 => X"7F10",
	216 => X"77AD",
	217 => X"6956",
	218 => X"54E0",
	219 => X"3B7B",
	220 => X"1EA1",
	221 => X"0000",
	222 => X"E15D",
	223 => X"C483",
	224 => X"AB1E",
	225 => X"96A8",
	226 => X"8851",
	227 => X"80EE",
	228 => X"80EE",
	229 => X"8851",
	230 => X"96A8",
	231 => X"AB1E",
	232 => X"C483",
	233 => X"E15D",
	234 => X"FFFE",
	235 => X"1EA1",
	236 => X"3B7B",
	237 => X"54E0",
	238 => X"6956",
	239 => X"77AD",
	240 => X"7F10",
	241 => X"7F10",
	242 => X"77AD",
	243 => X"6956",
	244 => X"54E0",
	245 => X"3B7B",
	246 => X"1EA1",
	247 => X"0000",
	others => X"0000"
);

BEGIN

--map all notes
key15_map: SampleContainer port map(clk, keys(15), C3, C4, C5, num_samples(015), num_samples(115), num_samples(215), octave, audio_request, k15);
key14_map: SampleContainer port map(clk, keys(14), CS3, CS4, CS5, num_samples(014), num_samples(114), num_samples(214), octave, audio_request, k14);
key13_map: SampleContainer port map(clk, keys(13), D3, D4, D5, num_samples(013), num_samples(113), num_samples(213), octave, audio_request, k13);
key12_map: SampleContainer port map(clk, keys(12), DS3, DS4, DS5, num_samples(012), num_samples(112), num_samples(212), octave, audio_request, k12);
key11_map: SampleContainer port map(clk, keys(11), E3, E4, E5, num_samples(011), num_samples(111), num_samples(211), octave, audio_request, k11);
key10_map: SampleContainer port map(clk, keys(10), F3, F4, F5, num_samples(010), num_samples(110), num_samples(210), octave, audio_request, k10);
key9_map: SampleContainer port map(clk, keys(9), FS3, FS4, FS5, num_samples(009), num_samples(109), num_samples(209), octave, audio_request, k9);
key8_map: SampleContainer port map(clk, keys(8), G3, G4, G5, num_samples(008), num_samples(108), num_samples(208), octave, audio_request, k8);
key7_map: SampleContainer port map(clk, keys(7), GS3, GS4, GS5, num_samples(007), num_samples(107), num_samples(207), octave, audio_request, k7);
key6_map: SampleContainer port map(clk, keys(6), A3, A4, A5, num_samples(006), num_samples(106), num_samples(206), octave, audio_request, k6);
key5_map: SampleContainer port map(clk, keys(5), AS3, AS4, AS5, num_samples(005), num_samples(105), num_samples(205), octave, audio_request, k5);
key4_map: SampleContainer port map(clk, keys(4), B3, B4, B5, num_samples(004), num_samples(104), num_samples(204), octave, audio_request, k4);
key3_map: SampleContainer port map(clk, keys(3), C4, C5, C6, num_samples(003), num_samples(103), num_samples(203), octave, audio_request, k3);
key2_map: SampleContainer port map(clk, keys(2), CS4, CS5, CS6, num_samples(002), num_samples(102), num_samples(202), octave, audio_request, k2);
key1_map: SampleContainer port map(clk, keys(1), D4, D5, D6, num_samples(001), num_samples(101), num_samples(201), octave, audio_request, k1);
key0_map: SampleContainer port map(clk, keys(0), DS4, DS5, DS6, num_samples(000), num_samples(100), num_samples(200), octave, audio_request, k0);

sample_adder: SampleAdder16 port map(keys, k0, k1, k2, k3, k4, k5, k6, k7, k8, k9, k10, k11, k12, k13, k14, k15, z);

END ARCHITECTURE rom;