library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.constants.all;

entity reverb is
	port(
		source_signal : in unsigned(DATA_SIZE - 1 downto 0);
		clear_bit, clk, switch: in std_logic;
		output: out unsigned(DATA_SIZE - 1 downto 0)
		);
end entity reverb;

architecture behavioral of reverb is

	component reverb_FIFO is
		generic(
			constant DATA_SIZE : positive := 16;
			constant FIFO_SIZE : positive := 48);
		port(
			clk : in std_logic;
			reset : in std_logic;
			write_enable : in std_logic;
			read_enable : in std_logic;
			data_in : in unsigned (DATA_SIZE - 1 downto 0);
			data_out : out unsigned (DATA_SIZE - 1 downto 0);
			empty : out std_logic;
			full : out std_logic);
	end component reverb_FIFO;
	
	component reverb_adder is
		port(
		IN1,IN2: in unsigned(DATA_SIZE - 1 downto 0);
		SUM    : out unsigned(DATA_SIZE - 1 downto 0));
	end component reverb_adder;
	
	component AND16 is
		port(
		A,B: in unsigned(DATA_SIZE - 1 downto 0);
		C  : out unsigned(DATA_SIZE - 1 downto 0));
	end component AND16;
	
	signal fifo_output, and_output: unsigned(DATA_SIZE - 1 downto 0);
	signal fifo_reset, fifo_write_en, fifo_read_en, fifo_empty, fifo_full : std_logic;
	signal fifo_in_data, fifo_out_data, AND_switch : unsigned (DATA_SIZE - 1 downto 0);
	
	begin
	
	FIFO_0: reverb_FIFO port map(clk, fifo_reset, fifo_write_en, fifo_read_en, fifo_in_data, fifo_out_data, fifo_empty, fifo_full);
	
	AND_0: AND16 port map(fifo_out_data, AND_switch, and_output);
	
	ADDER_0: reverb_adder port map(source_signal, and_output, output);
	
	process(switch) is begin
	if (switch = '0') then
	  AND_switch <= x"0000";
	else
	  AND_switch <= x"1111";
	end if;
	end process;
	  
	process(clk) is begin
	if (clear_bit = '1') then
	  fifo_reset <= '1';
	elsif(rising_edge(clk)) then
	  fifo_write_en <= '1';
	  fifo_read_en <= '1';
	end if;
	end process;

end behavioral;