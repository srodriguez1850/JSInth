library ieee;
use ieee.std_logic_1164.all;

package constants is
	constant DATA_SIZE : natural := 16;
	end package constants;
	
package body constants is
end package body constants;