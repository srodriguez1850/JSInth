LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE IEEE.std_logic_misc.all;
USE work.typeDeclarations.all;

ENTITY audioROM IS
PORT(
	clk: in std_logic;
	audio_request: in std_logic;
	keys: in std_logic_vector (15 downto 0);
	octave: in std_logic_vector (1 downto 0);
	z: out unsigned (15 downto 0)
);
END ENTITY audioROM;

ARCHITECTURE rom OF audioROM IS

COMPONENT SampleAdder16 IS
PORT(
		keys: in std_logic_vector(15 downto 0);

		a: in unsigned(15 downto 0);
		b: in unsigned(15 downto 0);
		c: in unsigned(15 downto 0);
		d: in unsigned(15 downto 0);
		e: in unsigned(15 downto 0);
		f: in unsigned(15 downto 0);
		g: in unsigned(15 downto 0);
		h: in unsigned(15 downto 0);
		i: in unsigned(15 downto 0);
		j: in unsigned(15 downto 0);
		k: in unsigned(15 downto 0);
		l: in unsigned(15 downto 0);
		m: in unsigned(15 downto 0);
		n: in unsigned(15 downto 0);
		o: in unsigned(15 downto 0);
		p: in unsigned(15 downto 0);
		
		z: out unsigned(15 downto 0)
);
END COMPONENT SampleAdder16;

COMPONENT SampleContainer IS
PORT(
		clk: in std_logic;
		stream: in std_logic;
		rom1, rom2, rom3: in hex;
		loop1, loop2, loop3: in natural;
		octave: in std_logic_vector (1 downto 0);
		audio_request: in std_logic;
		z: out unsigned (15 downto 0)
);
END COMPONENT SampleContainer;

SIGNAL k0, k1, k2, k3, k4, k5, k6, k7, k8, k9, k10, k11, k12, k13, k14, k15: unsigned (15 downto 0) := X"0000";

CONSTANT num_samples: nat_num := (
	--indexing set by octave(1) - tone(2)
	000 => 103,
	001 => 109,
	002 => 116,
	003 => 123,
	004 => 130,
	005 => 138,
	006 => 147,
	007 => 155,
	008 => 165,
	009 => 174,
	010 => 185,
	011 => 196,
	012 => 207,
	013 => 220,
	014 => 233,
	015 => 247,
	100 => 51,
	101 => 54,
	102 => 58,
	103 => 61,
	104 => 65,
	105 => 69,
	106 => 73,
	107 => 77,
	108 => 82,
	109 => 87,
	110 => 92,
	111 => 97,
	112 => 103,
	113 => 109,
	114 => 116,
	115 => 123,
	200 => 51,
	201 => 54,
	202 => 58,
	203 => 61,
	204 => 25,
	205 => 27,
	206 => 28,
	207 => 30,
	208 => 32,
	209 => 34,
	210 => 36,
	211 => 38,
	212 => 41,
	213 => 43,
	214 => 46,
	215 => 48,
	others => 0
);

CONSTANT C3: hex := (
	000 => X"0000",
	001 => X"033E",
	002 => X"067B",
	003 => X"09B8",
	004 => X"0CF2",
	005 => X"102B",
	006 => X"1361",
	007 => X"1694",
	008 => X"19C3",
	009 => X"1CEE",
	010 => X"2015",
	011 => X"2336",
	012 => X"2651",
	013 => X"2966",
	014 => X"2C74",
	015 => X"2F7A",
	016 => X"3279",
	017 => X"3570",
	018 => X"385E",
	019 => X"3B43",
	020 => X"3E1D",
	021 => X"40EE",
	022 => X"43B4",
	023 => X"466F",
	024 => X"491E",
	025 => X"4BC2",
	026 => X"4E58",
	027 => X"50E2",
	028 => X"535F",
	029 => X"55CE",
	030 => X"582F",
	031 => X"5A81",
	032 => X"5CC5",
	033 => X"5EF9",
	034 => X"611E",
	035 => X"6332",
	036 => X"6537",
	037 => X"672B",
	038 => X"690D",
	039 => X"6ADF",
	040 => X"6C9F",
	041 => X"6E4D",
	042 => X"6FE9",
	043 => X"7173",
	044 => X"72EA",
	045 => X"744E",
	046 => X"759F",
	047 => X"76DD",
	048 => X"7807",
	049 => X"791D",
	050 => X"7A20",
	051 => X"7B0E",
	052 => X"7BE8",
	053 => X"7CAE",
	054 => X"7D60",
	055 => X"7DFD",
	056 => X"7E85",
	057 => X"7EF8",
	058 => X"7F56",
	059 => X"7FA0",
	060 => X"7FD4",
	061 => X"7FF4",
	062 => X"7FFF",
	063 => X"7FF4",
	064 => X"7FD4",
	065 => X"7FA0",
	066 => X"7F56",
	067 => X"7EF8",
	068 => X"7E85",
	069 => X"7DFD",
	070 => X"7D60",
	071 => X"7CAE",
	072 => X"7BE8",
	073 => X"7B0E",
	074 => X"7A20",
	075 => X"791D",
	076 => X"7807",
	077 => X"76DD",
	078 => X"759F",
	079 => X"744E",
	080 => X"72EA",
	081 => X"7173",
	082 => X"6FE9",
	083 => X"6E4D",
	084 => X"6C9F",
	085 => X"6ADF",
	086 => X"690D",
	087 => X"672B",
	088 => X"6537",
	089 => X"6332",
	090 => X"611E",
	091 => X"5EF9",
	092 => X"5CC5",
	093 => X"5A81",
	094 => X"582F",
	095 => X"55CE",
	096 => X"535F",
	097 => X"50E2",
	098 => X"4E58",
	099 => X"4BC2",
	100 => X"491E",
	101 => X"466F",
	102 => X"43B4",
	103 => X"40EE",
	104 => X"3E1D",
	105 => X"3B43",
	106 => X"385E",
	107 => X"3570",
	108 => X"3279",
	109 => X"2F7A",
	110 => X"2C74",
	111 => X"2966",
	112 => X"2651",
	113 => X"2336",
	114 => X"2015",
	115 => X"1CEE",
	116 => X"19C3",
	117 => X"1694",
	118 => X"1361",
	119 => X"102B",
	120 => X"0CF2",
	121 => X"09B8",
	122 => X"067B",
	123 => X"033E",
	124 => X"0000",
	125 => X"FCBF",
	126 => X"F982",
	127 => X"F645",
	128 => X"F30B",
	129 => X"EFD2",
	130 => X"EC9C",
	131 => X"E969",
	132 => X"E63A",
	133 => X"E30F",
	134 => X"DFE8",
	135 => X"DCC7",
	136 => X"D9AC",
	137 => X"D697",
	138 => X"D389",
	139 => X"D083",
	140 => X"CD84",
	141 => X"CA8D",
	142 => X"C79F",
	143 => X"C4BA",
	144 => X"C1E0",
	145 => X"BF0F",
	146 => X"BC49",
	147 => X"B98E",
	148 => X"B6DF",
	149 => X"B43B",
	150 => X"B1A5",
	151 => X"AF1B",
	152 => X"AC9E",
	153 => X"AA2F",
	154 => X"A7CE",
	155 => X"A57C",
	156 => X"A338",
	157 => X"A104",
	158 => X"9EDF",
	159 => X"9CCB",
	160 => X"9AC6",
	161 => X"98D2",
	162 => X"96F0",
	163 => X"951E",
	164 => X"935E",
	165 => X"91B0",
	166 => X"9014",
	167 => X"8E8A",
	168 => X"8D13",
	169 => X"8BAF",
	170 => X"8A5E",
	171 => X"8920",
	172 => X"87F6",
	173 => X"86E0",
	174 => X"85DD",
	175 => X"84EF",
	176 => X"8415",
	177 => X"834F",
	178 => X"829D",
	179 => X"8200",
	180 => X"8178",
	181 => X"8105",
	182 => X"80A7",
	183 => X"805D",
	184 => X"8029",
	185 => X"8009",
	186 => X"7FFF",
	187 => X"8009",
	188 => X"8029",
	189 => X"805D",
	190 => X"80A7",
	191 => X"8105",
	192 => X"8178",
	193 => X"8200",
	194 => X"829D",
	195 => X"834F",
	196 => X"8415",
	197 => X"84EF",
	198 => X"85DD",
	199 => X"86E0",
	200 => X"87F6",
	201 => X"8920",
	202 => X"8A5E",
	203 => X"8BAF",
	204 => X"8D13",
	205 => X"8E8A",
	206 => X"9014",
	207 => X"91B0",
	208 => X"935E",
	209 => X"951E",
	210 => X"96F0",
	211 => X"98D2",
	212 => X"9AC6",
	213 => X"9CCB",
	214 => X"9EDF",
	215 => X"A104",
	216 => X"A338",
	217 => X"A57C",
	218 => X"A7CE",
	219 => X"AA2F",
	220 => X"AC9E",
	221 => X"AF1B",
	222 => X"B1A5",
	223 => X"B43B",
	224 => X"B6DF",
	225 => X"B98E",
	226 => X"BC49",
	227 => X"BF0F",
	228 => X"C1E0",
	229 => X"C4BA",
	230 => X"C79F",
	231 => X"CA8D",
	232 => X"CD84",
	233 => X"D083",
	234 => X"D389",
	235 => X"D697",
	236 => X"D9AC",
	237 => X"DCC7",
	238 => X"DFE8",
	239 => X"E30F",
	240 => X"E63A",
	241 => X"E969",
	242 => X"EC9C",
	243 => X"EFD2",
	244 => X"F30B",
	245 => X"F645",
	246 => X"F982",
	247 => X"FCBF",
	others => X"0000"
);

CONSTANT CS3: hex := (
	000 => X"0000",
	001 => X"036F",
	002 => X"06DE",
	003 => X"0A4C",
	004 => X"0DB8",
	005 => X"1121",
	006 => X"1488",
	007 => X"17EA",
	008 => X"1B48",
	009 => X"1EA1",
	010 => X"21F4",
	011 => X"2542",
	012 => X"2888",
	013 => X"2BC6",
	014 => X"2EFD",
	015 => X"322B",
	016 => X"3550",
	017 => X"386B",
	018 => X"3B7B",
	019 => X"3E81",
	020 => X"417A",
	021 => X"4468",
	022 => X"474A",
	023 => X"4A1E",
	024 => X"4CE4",
	025 => X"4F9C",
	026 => X"5246",
	027 => X"54E0",
	028 => X"576B",
	029 => X"59E5",
	030 => X"5C4F",
	031 => X"5EA8",
	032 => X"60EF",
	033 => X"6325",
	034 => X"6548",
	035 => X"6759",
	036 => X"6956",
	037 => X"6B40",
	038 => X"6D16",
	039 => X"6ED9",
	040 => X"7086",
	041 => X"721F",
	042 => X"73A3",
	043 => X"7511",
	044 => X"766A",
	045 => X"77AD",
	046 => X"78DA",
	047 => X"79F1",
	048 => X"7AF1",
	049 => X"7BDA",
	050 => X"7CAD",
	051 => X"7D68",
	052 => X"7E0D",
	053 => X"7E9A",
	054 => X"7F10",
	055 => X"7F6E",
	056 => X"7FB5",
	057 => X"7FE4",
	058 => X"7FFC",
	059 => X"7FFC",
	060 => X"7FE4",
	061 => X"7FB5",
	062 => X"7F6E",
	063 => X"7F10",
	064 => X"7E9A",
	065 => X"7E0D",
	066 => X"7D68",
	067 => X"7CAD",
	068 => X"7BDA",
	069 => X"7AF1",
	070 => X"79F1",
	071 => X"78DA",
	072 => X"77AD",
	073 => X"766A",
	074 => X"7511",
	075 => X"73A3",
	076 => X"721F",
	077 => X"7086",
	078 => X"6ED9",
	079 => X"6D16",
	080 => X"6B40",
	081 => X"6956",
	082 => X"6759",
	083 => X"6548",
	084 => X"6325",
	085 => X"60EF",
	086 => X"5EA8",
	087 => X"5C4F",
	088 => X"59E5",
	089 => X"576B",
	090 => X"54E0",
	091 => X"5246",
	092 => X"4F9C",
	093 => X"4CE4",
	094 => X"4A1E",
	095 => X"474A",
	096 => X"4468",
	097 => X"417A",
	098 => X"3E81",
	099 => X"3B7B",
	100 => X"386B",
	101 => X"3550",
	102 => X"322B",
	103 => X"2EFD",
	104 => X"2BC6",
	105 => X"2888",
	106 => X"2542",
	107 => X"21F4",
	108 => X"1EA1",
	109 => X"1B48",
	110 => X"17EA",
	111 => X"1488",
	112 => X"1121",
	113 => X"0DB8",
	114 => X"0A4C",
	115 => X"06DE",
	116 => X"036F",
	117 => X"FFFD",
	118 => X"FC8E",
	119 => X"F91F",
	120 => X"F5B1",
	121 => X"F245",
	122 => X"EEDC",
	123 => X"EB75",
	124 => X"E813",
	125 => X"E4B5",
	126 => X"E15C",
	127 => X"DE09",
	128 => X"DABB",
	129 => X"D775",
	130 => X"D437",
	131 => X"D100",
	132 => X"CDD2",
	133 => X"CAAD",
	134 => X"C792",
	135 => X"C482",
	136 => X"C17C",
	137 => X"BE83",
	138 => X"BB95",
	139 => X"B8B3",
	140 => X"B5DF",
	141 => X"B319",
	142 => X"B061",
	143 => X"ADB7",
	144 => X"AB1D",
	145 => X"A892",
	146 => X"A618",
	147 => X"A3AE",
	148 => X"A155",
	149 => X"9F0E",
	150 => X"9CD8",
	151 => X"9AB5",
	152 => X"98A4",
	153 => X"96A7",
	154 => X"94BD",
	155 => X"92E7",
	156 => X"9124",
	157 => X"8F77",
	158 => X"8DDE",
	159 => X"8C5A",
	160 => X"8AEC",
	161 => X"8993",
	162 => X"8850",
	163 => X"8723",
	164 => X"860C",
	165 => X"850C",
	166 => X"8423",
	167 => X"8350",
	168 => X"8295",
	169 => X"81F0",
	170 => X"8163",
	171 => X"80ED",
	172 => X"808F",
	173 => X"8048",
	174 => X"8019",
	175 => X"8001",
	176 => X"8001",
	177 => X"8019",
	178 => X"8048",
	179 => X"808F",
	180 => X"80ED",
	181 => X"8163",
	182 => X"81F0",
	183 => X"8295",
	184 => X"8350",
	185 => X"8423",
	186 => X"850C",
	187 => X"860C",
	188 => X"8723",
	189 => X"8850",
	190 => X"8993",
	191 => X"8AEC",
	192 => X"8C5A",
	193 => X"8DDE",
	194 => X"8F77",
	195 => X"9124",
	196 => X"92E7",
	197 => X"94BD",
	198 => X"96A7",
	199 => X"98A4",
	200 => X"9AB5",
	201 => X"9CD8",
	202 => X"9F0E",
	203 => X"A155",
	204 => X"A3AE",
	205 => X"A618",
	206 => X"A892",
	207 => X"AB1D",
	208 => X"ADB7",
	209 => X"B061",
	210 => X"B319",
	211 => X"B5DF",
	212 => X"B8B3",
	213 => X"BB95",
	214 => X"BE83",
	215 => X"C17C",
	216 => X"C482",
	217 => X"C792",
	218 => X"CAAD",
	219 => X"CDD2",
	220 => X"D100",
	221 => X"D437",
	222 => X"D775",
	223 => X"DABB",
	224 => X"DE09",
	225 => X"E15C",
	226 => X"E4B5",
	227 => X"E813",
	228 => X"EB75",
	229 => X"EEDC",
	230 => X"F245",
	231 => X"F5B1",
	232 => X"F91F",
	233 => X"FC8E",
	234 => X"0000",
	235 => X"036F",
	236 => X"06DE",
	237 => X"0A4C",
	238 => X"0DB8",
	239 => X"1121",
	240 => X"1488",
	241 => X"17EA",
	242 => X"1B48",
	243 => X"1EA1",
	244 => X"21F4",
	245 => X"2542",
	246 => X"2888",
	247 => X"2BC6",
	others => X"0000"
);

CONSTANT D3: hex := (
	000 => X"0000",
	001 => X"03A3",
	002 => X"0746",
	003 => X"0AE7",
	004 => X"0E86",
	005 => X"1222",
	006 => X"15BA",
	007 => X"194E",
	008 => X"1CDC",
	009 => X"2065",
	010 => X"23E6",
	011 => X"2761",
	012 => X"2AD3",
	013 => X"2E3C",
	014 => X"319C",
	015 => X"34F2",
	016 => X"383C",
	017 => X"3B7B",
	018 => X"3EAE",
	019 => X"41D3",
	020 => X"44EB",
	021 => X"47F5",
	022 => X"4AF0",
	023 => X"4DDB",
	024 => X"50B7",
	025 => X"5381",
	026 => X"563A",
	027 => X"58E2",
	028 => X"5B77",
	029 => X"5DF9",
	030 => X"6068",
	031 => X"62C2",
	032 => X"6509",
	033 => X"673A",
	034 => X"6956",
	035 => X"6B5C",
	036 => X"6D4C",
	037 => X"6F26",
	038 => X"70E8",
	039 => X"7293",
	040 => X"7427",
	041 => X"75A2",
	042 => X"7705",
	043 => X"784F",
	044 => X"7981",
	045 => X"7A99",
	046 => X"7B98",
	047 => X"7C7D",
	048 => X"7D49",
	049 => X"7DFB",
	050 => X"7E92",
	051 => X"7F10",
	052 => X"7F73",
	053 => X"7FBB",
	054 => X"7FEA",
	055 => X"7FFE",
	056 => X"7FF7",
	057 => X"7FD6",
	058 => X"7F9A",
	059 => X"7F44",
	060 => X"7ED4",
	061 => X"7E4A",
	062 => X"7DA5",
	063 => X"7CE6",
	064 => X"7C0E",
	065 => X"7B1C",
	066 => X"7A10",
	067 => X"78EB",
	068 => X"77AD",
	069 => X"7656",
	070 => X"74E7",
	071 => X"7360",
	072 => X"71C1",
	073 => X"700A",
	074 => X"6E3C",
	075 => X"6C57",
	076 => X"6A5C",
	077 => X"684B",
	078 => X"6624",
	079 => X"63E8",
	080 => X"6198",
	081 => X"5F33",
	082 => X"5CBA",
	083 => X"5A2F",
	084 => X"5790",
	085 => X"54E0",
	086 => X"521E",
	087 => X"4F4B",
	088 => X"4C68",
	089 => X"4974",
	090 => X"4672",
	091 => X"4361",
	092 => X"4042",
	093 => X"3D16",
	094 => X"39DD",
	095 => X"3698",
	096 => X"3348",
	097 => X"2FED",
	098 => X"2C89",
	099 => X"291B",
	100 => X"25A5",
	101 => X"2226",
	102 => X"1EA1",
	103 => X"1B16",
	104 => X"1784",
	105 => X"13EE",
	106 => X"1054",
	107 => X"0CB7",
	108 => X"0917",
	109 => X"0574",
	110 => X"01D1",
	111 => X"FE2C",
	112 => X"FA89",
	113 => X"F6E6",
	114 => X"F346",
	115 => X"EFA9",
	116 => X"EC0F",
	117 => X"E879",
	118 => X"E4E7",
	119 => X"E15C",
	120 => X"DDD7",
	121 => X"DA58",
	122 => X"D6E2",
	123 => X"D374",
	124 => X"D010",
	125 => X"CCB5",
	126 => X"C965",
	127 => X"C620",
	128 => X"C2E7",
	129 => X"BFBB",
	130 => X"BC9C",
	131 => X"B98B",
	132 => X"B689",
	133 => X"B395",
	134 => X"B0B2",
	135 => X"ADDF",
	136 => X"AB1D",
	137 => X"A86D",
	138 => X"A5CE",
	139 => X"A343",
	140 => X"A0CA",
	141 => X"9E65",
	142 => X"9C15",
	143 => X"99D9",
	144 => X"97B2",
	145 => X"95A1",
	146 => X"93A6",
	147 => X"91C1",
	148 => X"8FF3",
	149 => X"8E3C",
	150 => X"8C9D",
	151 => X"8B16",
	152 => X"89A7",
	153 => X"8850",
	154 => X"8712",
	155 => X"85ED",
	156 => X"84E1",
	157 => X"83EF",
	158 => X"8317",
	159 => X"8258",
	160 => X"81B3",
	161 => X"8129",
	162 => X"80B9",
	163 => X"8063",
	164 => X"8027",
	165 => X"8006",
	166 => X"7FFF",
	167 => X"8013",
	168 => X"8042",
	169 => X"808A",
	170 => X"80ED",
	171 => X"816B",
	172 => X"8202",
	173 => X"82B4",
	174 => X"8380",
	175 => X"8465",
	176 => X"8564",
	177 => X"867C",
	178 => X"87AE",
	179 => X"88F8",
	180 => X"8A5B",
	181 => X"8BD6",
	182 => X"8D6A",
	183 => X"8F15",
	184 => X"90D7",
	185 => X"92B1",
	186 => X"94A1",
	187 => X"96A7",
	188 => X"98C3",
	189 => X"9AF4",
	190 => X"9D3B",
	191 => X"9F95",
	192 => X"A204",
	193 => X"A486",
	194 => X"A71B",
	195 => X"A9C3",
	196 => X"AC7C",
	197 => X"AF46",
	198 => X"B222",
	199 => X"B50D",
	200 => X"B808",
	201 => X"BB12",
	202 => X"BE2A",
	203 => X"C14F",
	204 => X"C482",
	205 => X"C7C1",
	206 => X"CB0B",
	207 => X"CE61",
	208 => X"D1C1",
	209 => X"D52A",
	210 => X"D89C",
	211 => X"DC17",
	212 => X"DF98",
	213 => X"E321",
	214 => X"E6AF",
	215 => X"EA43",
	216 => X"EDDB",
	217 => X"F177",
	218 => X"F516",
	219 => X"F8B7",
	220 => X"FC5A",
	221 => X"0000",
	222 => X"03A3",
	223 => X"0746",
	224 => X"0AE7",
	225 => X"0E86",
	226 => X"1222",
	227 => X"15BA",
	228 => X"194E",
	229 => X"1CDC",
	230 => X"2065",
	231 => X"23E6",
	232 => X"2761",
	233 => X"2AD3",
	234 => X"2E3C",
	235 => X"319C",
	236 => X"34F2",
	237 => X"383C",
	238 => X"3B7B",
	239 => X"3EAE",
	240 => X"41D3",
	241 => X"44EB",
	242 => X"47F5",
	243 => X"4AF0",
	244 => X"4DDB",
	245 => X"50B7",
	246 => X"5381",
	247 => X"563A",
	others => X"0000"
);

CONSTANT DS3: hex := (
	000 => X"0000",
	001 => X"03DD",
	002 => X"07BA",
	003 => X"0B95",
	004 => X"0F6D",
	005 => X"1342",
	006 => X"1712",
	007 => X"1ADD",
	008 => X"1EA1",
	009 => X"225E",
	010 => X"2614",
	011 => X"29C0",
	012 => X"2D63",
	013 => X"30FB",
	014 => X"3487",
	015 => X"3808",
	016 => X"3B7B",
	017 => X"3EE0",
	018 => X"4237",
	019 => X"457E",
	020 => X"48B5",
	021 => X"4BDB",
	022 => X"4EF0",
	023 => X"51F1",
	024 => X"54E0",
	025 => X"57BB",
	026 => X"5A81",
	027 => X"5D32",
	028 => X"5FCE",
	029 => X"6253",
	030 => X"64C1",
	031 => X"6718",
	032 => X"6956",
	033 => X"6B7C",
	034 => X"6D89",
	035 => X"6F7C",
	036 => X"7155",
	037 => X"7314",
	038 => X"74B8",
	039 => X"7640",
	040 => X"77AD",
	041 => X"78FE",
	042 => X"7A33",
	043 => X"7B4B",
	044 => X"7C46",
	045 => X"7D25",
	046 => X"7DE6",
	047 => X"7E89",
	048 => X"7F10",
	049 => X"7F78",
	050 => X"7FC3",
	051 => X"7FF0",
	052 => X"7FFF",
	053 => X"7FF0",
	054 => X"7FC3",
	055 => X"7F78",
	056 => X"7F10",
	057 => X"7E89",
	058 => X"7DE6",
	059 => X"7D25",
	060 => X"7C46",
	061 => X"7B4B",
	062 => X"7A33",
	063 => X"78FE",
	064 => X"77AD",
	065 => X"7640",
	066 => X"74B8",
	067 => X"7314",
	068 => X"7155",
	069 => X"6F7C",
	070 => X"6D89",
	071 => X"6B7C",
	072 => X"6956",
	073 => X"6718",
	074 => X"64C1",
	075 => X"6253",
	076 => X"5FCE",
	077 => X"5D32",
	078 => X"5A81",
	079 => X"57BB",
	080 => X"54E0",
	081 => X"51F1",
	082 => X"4EF0",
	083 => X"4BDB",
	084 => X"48B5",
	085 => X"457E",
	086 => X"4237",
	087 => X"3EE0",
	088 => X"3B7B",
	089 => X"3808",
	090 => X"3487",
	091 => X"30FB",
	092 => X"2D63",
	093 => X"29C0",
	094 => X"2614",
	095 => X"225E",
	096 => X"1EA1",
	097 => X"1ADD",
	098 => X"1712",
	099 => X"1342",
	100 => X"0F6D",
	101 => X"0B95",
	102 => X"07BA",
	103 => X"03DD",
	104 => X"0000",
	105 => X"FC20",
	106 => X"F843",
	107 => X"F468",
	108 => X"F090",
	109 => X"ECBB",
	110 => X"E8EB",
	111 => X"E520",
	112 => X"E15C",
	113 => X"DD9F",
	114 => X"D9E9",
	115 => X"D63D",
	116 => X"D29A",
	117 => X"CF02",
	118 => X"CB76",
	119 => X"C7F5",
	120 => X"C482",
	121 => X"C11D",
	122 => X"BDC6",
	123 => X"BA7F",
	124 => X"B748",
	125 => X"B422",
	126 => X"B10D",
	127 => X"AE0C",
	128 => X"AB1D",
	129 => X"A842",
	130 => X"A57C",
	131 => X"A2CB",
	132 => X"A02F",
	133 => X"9DAA",
	134 => X"9B3C",
	135 => X"98E5",
	136 => X"96A7",
	137 => X"9481",
	138 => X"9274",
	139 => X"9081",
	140 => X"8EA8",
	141 => X"8CE9",
	142 => X"8B45",
	143 => X"89BD",
	144 => X"8850",
	145 => X"86FF",
	146 => X"85CA",
	147 => X"84B2",
	148 => X"83B7",
	149 => X"82D8",
	150 => X"8217",
	151 => X"8174",
	152 => X"80ED",
	153 => X"8085",
	154 => X"803A",
	155 => X"800D",
	156 => X"7FFF",
	157 => X"800D",
	158 => X"803A",
	159 => X"8085",
	160 => X"80ED",
	161 => X"8174",
	162 => X"8217",
	163 => X"82D8",
	164 => X"83B7",
	165 => X"84B2",
	166 => X"85CA",
	167 => X"86FF",
	168 => X"8850",
	169 => X"89BD",
	170 => X"8B45",
	171 => X"8CE9",
	172 => X"8EA8",
	173 => X"9081",
	174 => X"9274",
	175 => X"9481",
	176 => X"96A7",
	177 => X"98E5",
	178 => X"9B3C",
	179 => X"9DAA",
	180 => X"A02F",
	181 => X"A2CB",
	182 => X"A57C",
	183 => X"A842",
	184 => X"AB1D",
	185 => X"AE0C",
	186 => X"B10D",
	187 => X"B422",
	188 => X"B748",
	189 => X"BA7F",
	190 => X"BDC6",
	191 => X"C11D",
	192 => X"C482",
	193 => X"C7F5",
	194 => X"CB76",
	195 => X"CF02",
	196 => X"D29A",
	197 => X"D63D",
	198 => X"D9E9",
	199 => X"DD9F",
	200 => X"E15C",
	201 => X"E520",
	202 => X"E8EB",
	203 => X"ECBB",
	204 => X"F090",
	205 => X"F468",
	206 => X"F843",
	207 => X"FC20",
	208 => X"FFFD",
	209 => X"03DD",
	210 => X"07BA",
	211 => X"0B95",
	212 => X"0F6D",
	213 => X"1342",
	214 => X"1712",
	215 => X"1ADD",
	216 => X"1EA1",
	217 => X"225E",
	218 => X"2614",
	219 => X"29C0",
	220 => X"2D63",
	221 => X"30FB",
	222 => X"3487",
	223 => X"3808",
	224 => X"3B7B",
	225 => X"3EE0",
	226 => X"4237",
	227 => X"457E",
	228 => X"48B5",
	229 => X"4BDB",
	230 => X"4EF0",
	231 => X"51F1",
	232 => X"54E0",
	233 => X"57BB",
	234 => X"5A81",
	235 => X"5D32",
	236 => X"5FCE",
	237 => X"6253",
	238 => X"64C1",
	239 => X"6718",
	240 => X"6956",
	241 => X"6B7C",
	242 => X"6D89",
	243 => X"6F7C",
	244 => X"7155",
	245 => X"7314",
	246 => X"74B8",
	247 => X"7640",
	others => X"0000"
);

CONSTANT E3: hex := (
	000 => X"0000",
	001 => X"0414",
	002 => X"0828",
	003 => X"0C3A",
	004 => X"1048",
	005 => X"1453",
	006 => X"1858",
	007 => X"1C56",
	008 => X"204E",
	009 => X"243D",
	010 => X"2822",
	011 => X"2BFD",
	012 => X"2FCD",
	013 => X"3390",
	014 => X"3745",
	015 => X"3AED",
	016 => X"3E84",
	017 => X"420C",
	018 => X"4583",
	019 => X"48E7",
	020 => X"4C38",
	021 => X"4F76",
	022 => X"529F",
	023 => X"55B2",
	024 => X"58AF",
	025 => X"5B95",
	026 => X"5E63",
	027 => X"6118",
	028 => X"63B4",
	029 => X"6637",
	030 => X"689E",
	031 => X"6AEB",
	032 => X"6D1B",
	033 => X"6F2F",
	034 => X"7126",
	035 => X"7300",
	036 => X"74BC",
	037 => X"7659",
	038 => X"77D8",
	039 => X"7937",
	040 => X"7A77",
	041 => X"7B97",
	042 => X"7C96",
	043 => X"7D76",
	044 => X"7E34",
	045 => X"7ED2",
	046 => X"7F4F",
	047 => X"7FAA",
	048 => X"7FE4",
	049 => X"7FFD",
	050 => X"7FF5",
	051 => X"7FCB",
	052 => X"7F81",
	053 => X"7F14",
	054 => X"7E87",
	055 => X"7DD9",
	056 => X"7D0A",
	057 => X"7C1B",
	058 => X"7B0B",
	059 => X"79DB",
	060 => X"788B",
	061 => X"771C",
	062 => X"758E",
	063 => X"73E2",
	064 => X"7217",
	065 => X"702E",
	066 => X"6E29",
	067 => X"6C06",
	068 => X"69C8",
	069 => X"676E",
	070 => X"64F9",
	071 => X"626A",
	072 => X"5FC1",
	073 => X"5CFF",
	074 => X"5A25",
	075 => X"5733",
	076 => X"542B",
	077 => X"510D",
	078 => X"4DDA",
	079 => X"4A92",
	080 => X"4737",
	081 => X"43CA",
	082 => X"404A",
	083 => X"3CBA",
	084 => X"391B",
	085 => X"356C",
	086 => X"31B0",
	087 => X"2DE6",
	088 => X"2A11",
	089 => X"2631",
	090 => X"2246",
	091 => X"1E53",
	092 => X"1A58",
	093 => X"1656",
	094 => X"124E",
	095 => X"0E42",
	096 => X"0A31",
	097 => X"061F",
	098 => X"020A",
	099 => X"FDF3",
	100 => X"F9DE",
	101 => X"F5CC",
	102 => X"F1BB",
	103 => X"EDAF",
	104 => X"E9A7",
	105 => X"E5A5",
	106 => X"E1AA",
	107 => X"DDB7",
	108 => X"D9CC",
	109 => X"D5EC",
	110 => X"D217",
	111 => X"CE4D",
	112 => X"CA91",
	113 => X"C6E2",
	114 => X"C343",
	115 => X"BFB3",
	116 => X"BC33",
	117 => X"B8C6",
	118 => X"B56B",
	119 => X"B223",
	120 => X"AEF0",
	121 => X"ABD2",
	122 => X"A8CA",
	123 => X"A5D8",
	124 => X"A2FE",
	125 => X"A03C",
	126 => X"9D93",
	127 => X"9B04",
	128 => X"988F",
	129 => X"9635",
	130 => X"93F7",
	131 => X"91D4",
	132 => X"8FCF",
	133 => X"8DE6",
	134 => X"8C1B",
	135 => X"8A6F",
	136 => X"88E1",
	137 => X"8772",
	138 => X"8622",
	139 => X"84F2",
	140 => X"83E2",
	141 => X"82F3",
	142 => X"8224",
	143 => X"8176",
	144 => X"80E9",
	145 => X"807C",
	146 => X"8032",
	147 => X"8008",
	148 => X"8000",
	149 => X"8019",
	150 => X"8053",
	151 => X"80AE",
	152 => X"812B",
	153 => X"81C9",
	154 => X"8287",
	155 => X"8367",
	156 => X"8466",
	157 => X"8586",
	158 => X"86C6",
	159 => X"8825",
	160 => X"89A4",
	161 => X"8B41",
	162 => X"8CFD",
	163 => X"8ED7",
	164 => X"90CE",
	165 => X"92E2",
	166 => X"9512",
	167 => X"975F",
	168 => X"99C6",
	169 => X"9C49",
	170 => X"9EE5",
	171 => X"A19A",
	172 => X"A468",
	173 => X"A74E",
	174 => X"AA4B",
	175 => X"AD5E",
	176 => X"B087",
	177 => X"B3C5",
	178 => X"B716",
	179 => X"BA7A",
	180 => X"BDF1",
	181 => X"C179",
	182 => X"C510",
	183 => X"C8B8",
	184 => X"CC6D",
	185 => X"D030",
	186 => X"D400",
	187 => X"D7DB",
	188 => X"DBC0",
	189 => X"DFAF",
	190 => X"E3A7",
	191 => X"E7A5",
	192 => X"EBAA",
	193 => X"EFB5",
	194 => X"F3C3",
	195 => X"F7D5",
	196 => X"FBE9",
	197 => X"0000",
	198 => X"0414",
	199 => X"0828",
	200 => X"0C3A",
	201 => X"1048",
	202 => X"1453",
	203 => X"1858",
	204 => X"1C56",
	205 => X"204E",
	206 => X"243D",
	207 => X"2822",
	208 => X"2BFD",
	209 => X"2FCD",
	210 => X"3390",
	211 => X"3745",
	212 => X"3AED",
	213 => X"3E84",
	214 => X"420C",
	215 => X"4583",
	216 => X"48E7",
	217 => X"4C38",
	218 => X"4F76",
	219 => X"529F",
	220 => X"55B2",
	221 => X"58AF",
	222 => X"5B95",
	223 => X"5E63",
	224 => X"6118",
	225 => X"63B4",
	226 => X"6637",
	227 => X"689E",
	228 => X"6AEB",
	229 => X"6D1B",
	230 => X"6F2F",
	231 => X"7126",
	232 => X"7300",
	233 => X"74BC",
	234 => X"7659",
	235 => X"77D8",
	236 => X"7937",
	237 => X"7A77",
	238 => X"7B97",
	239 => X"7C96",
	240 => X"7D76",
	241 => X"7E34",
	242 => X"7ED2",
	243 => X"7F4F",
	244 => X"7FAA",
	245 => X"7FE4",
	246 => X"7FFD",
	247 => X"7FF5",
	others => X"0000"
);

CONSTANT F3: hex := (
	000 => X"0000",
	001 => X"0452",
	002 => X"08A4",
	003 => X"0CF2",
	004 => X"113E",
	005 => X"1584",
	006 => X"19C3",
	007 => X"1DFC",
	008 => X"222B",
	009 => X"2651",
	010 => X"2A6B",
	011 => X"2E79",
	012 => X"3279",
	013 => X"366B",
	014 => X"3A4D",
	015 => X"3E1D",
	016 => X"41DC",
	017 => X"4587",
	018 => X"491E",
	019 => X"4CA0",
	020 => X"500B",
	021 => X"535F",
	022 => X"569B",
	023 => X"59BD",
	024 => X"5CC5",
	025 => X"5FB2",
	026 => X"6283",
	027 => X"6537",
	028 => X"67CD",
	029 => X"6A46",
	030 => X"6C9F",
	031 => X"6ED9",
	032 => X"70F2",
	033 => X"72EA",
	034 => X"74C0",
	035 => X"7675",
	036 => X"7807",
	037 => X"7976",
	038 => X"7AC1",
	039 => X"7BE8",
	040 => X"7CEC",
	041 => X"7DCB",
	042 => X"7E85",
	043 => X"7F1A",
	044 => X"7F8A",
	045 => X"7FD4",
	046 => X"7FFA",
	047 => X"7FFA",
	048 => X"7FD4",
	049 => X"7F8A",
	050 => X"7F1A",
	051 => X"7E85",
	052 => X"7DCB",
	053 => X"7CEC",
	054 => X"7BE8",
	055 => X"7AC1",
	056 => X"7976",
	057 => X"7807",
	058 => X"7675",
	059 => X"74C0",
	060 => X"72EA",
	061 => X"70F2",
	062 => X"6ED9",
	063 => X"6C9F",
	064 => X"6A46",
	065 => X"67CD",
	066 => X"6537",
	067 => X"6283",
	068 => X"5FB2",
	069 => X"5CC5",
	070 => X"59BD",
	071 => X"569B",
	072 => X"535F",
	073 => X"500B",
	074 => X"4CA0",
	075 => X"491E",
	076 => X"4587",
	077 => X"41DC",
	078 => X"3E1D",
	079 => X"3A4D",
	080 => X"366B",
	081 => X"3279",
	082 => X"2E79",
	083 => X"2A6B",
	084 => X"2651",
	085 => X"222B",
	086 => X"1DFC",
	087 => X"19C3",
	088 => X"1584",
	089 => X"113E",
	090 => X"0CF2",
	091 => X"08A4",
	092 => X"0452",
	093 => X"FFFD",
	094 => X"FBAB",
	095 => X"F759",
	096 => X"F30B",
	097 => X"EEBF",
	098 => X"EA79",
	099 => X"E63A",
	100 => X"E201",
	101 => X"DDD2",
	102 => X"D9AC",
	103 => X"D592",
	104 => X"D184",
	105 => X"CD84",
	106 => X"C992",
	107 => X"C5B0",
	108 => X"C1E0",
	109 => X"BE21",
	110 => X"BA76",
	111 => X"B6DF",
	112 => X"B35D",
	113 => X"AFF2",
	114 => X"AC9E",
	115 => X"A962",
	116 => X"A640",
	117 => X"A338",
	118 => X"A04B",
	119 => X"9D7A",
	120 => X"9AC6",
	121 => X"9830",
	122 => X"95B7",
	123 => X"935E",
	124 => X"9124",
	125 => X"8F0B",
	126 => X"8D13",
	127 => X"8B3D",
	128 => X"8988",
	129 => X"87F6",
	130 => X"8687",
	131 => X"853C",
	132 => X"8415",
	133 => X"8311",
	134 => X"8232",
	135 => X"8178",
	136 => X"80E3",
	137 => X"8073",
	138 => X"8029",
	139 => X"8003",
	140 => X"8003",
	141 => X"8029",
	142 => X"8073",
	143 => X"80E3",
	144 => X"8178",
	145 => X"8232",
	146 => X"8311",
	147 => X"8415",
	148 => X"853C",
	149 => X"8687",
	150 => X"87F6",
	151 => X"8988",
	152 => X"8B3D",
	153 => X"8D13",
	154 => X"8F0B",
	155 => X"9124",
	156 => X"935E",
	157 => X"95B7",
	158 => X"9830",
	159 => X"9AC6",
	160 => X"9D7A",
	161 => X"A04B",
	162 => X"A338",
	163 => X"A640",
	164 => X"A962",
	165 => X"AC9E",
	166 => X"AFF2",
	167 => X"B35D",
	168 => X"B6DF",
	169 => X"BA76",
	170 => X"BE21",
	171 => X"C1E0",
	172 => X"C5B0",
	173 => X"C992",
	174 => X"CD84",
	175 => X"D184",
	176 => X"D592",
	177 => X"D9AC",
	178 => X"DDD2",
	179 => X"E201",
	180 => X"E63A",
	181 => X"EA79",
	182 => X"EEBF",
	183 => X"F30B",
	184 => X"F759",
	185 => X"FBAB",
	186 => X"0000",
	187 => X"0452",
	188 => X"08A4",
	189 => X"0CF2",
	190 => X"113E",
	191 => X"1584",
	192 => X"19C3",
	193 => X"1DFC",
	194 => X"222B",
	195 => X"2651",
	196 => X"2A6B",
	197 => X"2E79",
	198 => X"3279",
	199 => X"366B",
	200 => X"3A4D",
	201 => X"3E1D",
	202 => X"41DC",
	203 => X"4587",
	204 => X"491E",
	205 => X"4CA0",
	206 => X"500B",
	207 => X"535F",
	208 => X"569B",
	209 => X"59BD",
	210 => X"5CC5",
	211 => X"5FB2",
	212 => X"6283",
	213 => X"6537",
	214 => X"67CD",
	215 => X"6A46",
	216 => X"6C9F",
	217 => X"6ED9",
	218 => X"70F2",
	219 => X"72EA",
	220 => X"74C0",
	221 => X"7675",
	222 => X"7807",
	223 => X"7976",
	224 => X"7AC1",
	225 => X"7BE8",
	226 => X"7CEC",
	227 => X"7DCB",
	228 => X"7E85",
	229 => X"7F1A",
	230 => X"7F8A",
	231 => X"7FD4",
	232 => X"7FFA",
	233 => X"7FFA",
	234 => X"7FD4",
	235 => X"7F8A",
	236 => X"7F1A",
	237 => X"7E85",
	238 => X"7DCB",
	239 => X"7CEC",
	240 => X"7BE8",
	241 => X"7AC1",
	242 => X"7976",
	243 => X"7807",
	244 => X"7675",
	245 => X"74C0",
	246 => X"72EA",
	247 => X"70F2",
	others => X"0000"
);

CONSTANT FS3: hex := (
	000 => X"0000",
	001 => X"0498",
	002 => X"092E",
	003 => X"0DC2",
	004 => X"1251",
	005 => X"16DA",
	006 => X"1B5C",
	007 => X"1FD4",
	008 => X"2442",
	009 => X"28A4",
	010 => X"2CF9",
	011 => X"313F",
	012 => X"3574",
	013 => X"3998",
	014 => X"3DA9",
	015 => X"41A6",
	016 => X"458D",
	017 => X"495C",
	018 => X"4D14",
	019 => X"50B3",
	020 => X"5436",
	021 => X"579E",
	022 => X"5AE9",
	023 => X"5E16",
	024 => X"6124",
	025 => X"6412",
	026 => X"66DF",
	027 => X"698A",
	028 => X"6C12",
	029 => X"6E76",
	030 => X"70B6",
	031 => X"72D1",
	032 => X"74C6",
	033 => X"7694",
	034 => X"783B",
	035 => X"79BB",
	036 => X"7B12",
	037 => X"7C41",
	038 => X"7D47",
	039 => X"7E23",
	040 => X"7ED6",
	041 => X"7F5F",
	042 => X"7FBE",
	043 => X"7FF3",
	044 => X"7FFD",
	045 => X"7FDE",
	046 => X"7F94",
	047 => X"7F20",
	048 => X"7E82",
	049 => X"7DBA",
	050 => X"7CC9",
	051 => X"7BAF",
	052 => X"7A6C",
	053 => X"7900",
	054 => X"776D",
	055 => X"75B2",
	056 => X"73D0",
	057 => X"71C8",
	058 => X"6F9B",
	059 => X"6D48",
	060 => X"6AD2",
	061 => X"6838",
	062 => X"657C",
	063 => X"629F",
	064 => X"5FA1",
	065 => X"5C83",
	066 => X"5947",
	067 => X"55EE",
	068 => X"5278",
	069 => X"4EE7",
	070 => X"4B3B",
	071 => X"4777",
	072 => X"439C",
	073 => X"3FAA",
	074 => X"3BA3",
	075 => X"3789",
	076 => X"335C",
	077 => X"2F1E",
	078 => X"2AD0",
	079 => X"2675",
	080 => X"220D",
	081 => X"1D99",
	082 => X"191C",
	083 => X"1497",
	084 => X"100A",
	085 => X"0B79",
	086 => X"06E3",
	087 => X"024C",
	088 => X"FDB1",
	089 => X"F91A",
	090 => X"F484",
	091 => X"EFF3",
	092 => X"EB66",
	093 => X"E6E1",
	094 => X"E264",
	095 => X"DDF0",
	096 => X"D988",
	097 => X"D52D",
	098 => X"D0DF",
	099 => X"CCA1",
	100 => X"C874",
	101 => X"C45A",
	102 => X"C053",
	103 => X"BC61",
	104 => X"B886",
	105 => X"B4C2",
	106 => X"B116",
	107 => X"AD85",
	108 => X"AA0F",
	109 => X"A6B6",
	110 => X"A37A",
	111 => X"A05C",
	112 => X"9D5E",
	113 => X"9A81",
	114 => X"97C5",
	115 => X"952B",
	116 => X"92B5",
	117 => X"9062",
	118 => X"8E35",
	119 => X"8C2D",
	120 => X"8A4B",
	121 => X"8890",
	122 => X"86FD",
	123 => X"8591",
	124 => X"844E",
	125 => X"8334",
	126 => X"8243",
	127 => X"817B",
	128 => X"80DD",
	129 => X"8069",
	130 => X"801F",
	131 => X"8000",
	132 => X"800A",
	133 => X"803F",
	134 => X"809E",
	135 => X"8127",
	136 => X"81DA",
	137 => X"82B6",
	138 => X"83BC",
	139 => X"84EB",
	140 => X"8642",
	141 => X"87C2",
	142 => X"8969",
	143 => X"8B37",
	144 => X"8D2C",
	145 => X"8F47",
	146 => X"9187",
	147 => X"93EB",
	148 => X"9673",
	149 => X"991E",
	150 => X"9BEB",
	151 => X"9ED9",
	152 => X"A1E7",
	153 => X"A514",
	154 => X"A85F",
	155 => X"ABC7",
	156 => X"AF4A",
	157 => X"B2E9",
	158 => X"B6A1",
	159 => X"BA70",
	160 => X"BE57",
	161 => X"C254",
	162 => X"C665",
	163 => X"CA89",
	164 => X"CEBE",
	165 => X"D304",
	166 => X"D759",
	167 => X"DBBB",
	168 => X"E029",
	169 => X"E4A1",
	170 => X"E923",
	171 => X"EDAC",
	172 => X"F23B",
	173 => X"F6CF",
	174 => X"FB65",
	175 => X"0000",
	176 => X"0498",
	177 => X"092E",
	178 => X"0DC2",
	179 => X"1251",
	180 => X"16DA",
	181 => X"1B5C",
	182 => X"1FD4",
	183 => X"2442",
	184 => X"28A4",
	185 => X"2CF9",
	186 => X"313F",
	187 => X"3574",
	188 => X"3998",
	189 => X"3DA9",
	190 => X"41A6",
	191 => X"458D",
	192 => X"495C",
	193 => X"4D14",
	194 => X"50B3",
	195 => X"5436",
	196 => X"579E",
	197 => X"5AE9",
	198 => X"5E16",
	199 => X"6124",
	200 => X"6412",
	201 => X"66DF",
	202 => X"698A",
	203 => X"6C12",
	204 => X"6E76",
	205 => X"70B6",
	206 => X"72D1",
	207 => X"74C6",
	208 => X"7694",
	209 => X"783B",
	210 => X"79BB",
	211 => X"7B12",
	212 => X"7C41",
	213 => X"7D47",
	214 => X"7E23",
	215 => X"7ED6",
	216 => X"7F5F",
	217 => X"7FBE",
	218 => X"7FF3",
	219 => X"7FFD",
	220 => X"7FDE",
	221 => X"7F94",
	222 => X"7F20",
	223 => X"7E82",
	224 => X"7DBA",
	225 => X"7CC9",
	226 => X"7BAF",
	227 => X"7A6C",
	228 => X"7900",
	229 => X"776D",
	230 => X"75B2",
	231 => X"73D0",
	232 => X"71C8",
	233 => X"6F9B",
	234 => X"6D48",
	235 => X"6AD2",
	236 => X"6838",
	237 => X"657C",
	238 => X"629F",
	239 => X"5FA1",
	240 => X"5C83",
	241 => X"5947",
	242 => X"55EE",
	243 => X"5278",
	244 => X"4EE7",
	245 => X"4B3B",
	246 => X"4777",
	247 => X"439C",
	others => X"0000"
);

CONSTANT G3: hex := (
	000 => X"0000",
	001 => X"04D7",
	002 => X"09AE",
	003 => X"0E80",
	004 => X"134E",
	005 => X"1814",
	006 => X"1CD1",
	007 => X"2184",
	008 => X"262B",
	009 => X"2AC3",
	010 => X"2F4C",
	011 => X"33C3",
	012 => X"3828",
	013 => X"3C78",
	014 => X"40B2",
	015 => X"44D4",
	016 => X"48DD",
	017 => X"4CCB",
	018 => X"509D",
	019 => X"5451",
	020 => X"57E6",
	021 => X"5B5B",
	022 => X"5EAF",
	023 => X"61E0",
	024 => X"64ED",
	025 => X"67D5",
	026 => X"6A97",
	027 => X"6D32",
	028 => X"6FA5",
	029 => X"71EF",
	030 => X"740F",
	031 => X"7605",
	032 => X"77CF",
	033 => X"796D",
	034 => X"7ADF",
	035 => X"7C24",
	036 => X"7D3B",
	037 => X"7E24",
	038 => X"7EDF",
	039 => X"7F6C",
	040 => X"7FCA",
	041 => X"7FF9",
	042 => X"7FF9",
	043 => X"7FCA",
	044 => X"7F6C",
	045 => X"7EDF",
	046 => X"7E24",
	047 => X"7D3B",
	048 => X"7C24",
	049 => X"7ADF",
	050 => X"796D",
	051 => X"77CF",
	052 => X"7605",
	053 => X"740F",
	054 => X"71EF",
	055 => X"6FA5",
	056 => X"6D32",
	057 => X"6A97",
	058 => X"67D5",
	059 => X"64ED",
	060 => X"61E0",
	061 => X"5EAF",
	062 => X"5B5B",
	063 => X"57E6",
	064 => X"5451",
	065 => X"509D",
	066 => X"4CCB",
	067 => X"48DD",
	068 => X"44D4",
	069 => X"40B2",
	070 => X"3C78",
	071 => X"3828",
	072 => X"33C3",
	073 => X"2F4C",
	074 => X"2AC3",
	075 => X"262B",
	076 => X"2184",
	077 => X"1CD1",
	078 => X"1814",
	079 => X"134E",
	080 => X"0E80",
	081 => X"09AE",
	082 => X"04D7",
	083 => X"0000",
	084 => X"FB26",
	085 => X"F64F",
	086 => X"F17D",
	087 => X"ECAF",
	088 => X"E7E9",
	089 => X"E32C",
	090 => X"DE79",
	091 => X"D9D2",
	092 => X"D53A",
	093 => X"D0B1",
	094 => X"CC3A",
	095 => X"C7D5",
	096 => X"C385",
	097 => X"BF4B",
	098 => X"BB29",
	099 => X"B720",
	100 => X"B332",
	101 => X"AF60",
	102 => X"ABAC",
	103 => X"A817",
	104 => X"A4A2",
	105 => X"A14E",
	106 => X"9E1D",
	107 => X"9B10",
	108 => X"9828",
	109 => X"9566",
	110 => X"92CB",
	111 => X"9058",
	112 => X"8E0E",
	113 => X"8BEE",
	114 => X"89F8",
	115 => X"882E",
	116 => X"8690",
	117 => X"851E",
	118 => X"83D9",
	119 => X"82C2",
	120 => X"81D9",
	121 => X"811E",
	122 => X"8091",
	123 => X"8033",
	124 => X"8004",
	125 => X"8004",
	126 => X"8033",
	127 => X"8091",
	128 => X"811E",
	129 => X"81D9",
	130 => X"82C2",
	131 => X"83D9",
	132 => X"851E",
	133 => X"8690",
	134 => X"882E",
	135 => X"89F8",
	136 => X"8BEE",
	137 => X"8E0E",
	138 => X"9058",
	139 => X"92CB",
	140 => X"9566",
	141 => X"9828",
	142 => X"9B10",
	143 => X"9E1D",
	144 => X"A14E",
	145 => X"A4A2",
	146 => X"A817",
	147 => X"ABAC",
	148 => X"AF60",
	149 => X"B332",
	150 => X"B720",
	151 => X"BB29",
	152 => X"BF4B",
	153 => X"C385",
	154 => X"C7D5",
	155 => X"CC3A",
	156 => X"D0B1",
	157 => X"D53A",
	158 => X"D9D2",
	159 => X"DE79",
	160 => X"E32C",
	161 => X"E7E9",
	162 => X"ECAF",
	163 => X"F17D",
	164 => X"F64F",
	165 => X"FB26",
	166 => X"0000",
	167 => X"04D7",
	168 => X"09AE",
	169 => X"0E80",
	170 => X"134E",
	171 => X"1814",
	172 => X"1CD1",
	173 => X"2184",
	174 => X"262B",
	175 => X"2AC3",
	176 => X"2F4C",
	177 => X"33C3",
	178 => X"3828",
	179 => X"3C78",
	180 => X"40B2",
	181 => X"44D4",
	182 => X"48DD",
	183 => X"4CCB",
	184 => X"509D",
	185 => X"5451",
	186 => X"57E6",
	187 => X"5B5B",
	188 => X"5EAF",
	189 => X"61E0",
	190 => X"64ED",
	191 => X"67D5",
	192 => X"6A97",
	193 => X"6D32",
	194 => X"6FA5",
	195 => X"71EF",
	196 => X"740F",
	197 => X"7605",
	198 => X"77CF",
	199 => X"796D",
	200 => X"7ADF",
	201 => X"7C24",
	202 => X"7D3B",
	203 => X"7E24",
	204 => X"7EDF",
	205 => X"7F6C",
	206 => X"7FCA",
	207 => X"7FF9",
	208 => X"7FF9",
	209 => X"7FCA",
	210 => X"7F6C",
	211 => X"7EDF",
	212 => X"7E24",
	213 => X"7D3B",
	214 => X"7C24",
	215 => X"7ADF",
	216 => X"796D",
	217 => X"77CF",
	218 => X"7605",
	219 => X"740F",
	220 => X"71EF",
	221 => X"6FA5",
	222 => X"6D32",
	223 => X"6A97",
	224 => X"67D5",
	225 => X"64ED",
	226 => X"61E0",
	227 => X"5EAF",
	228 => X"5B5B",
	229 => X"57E6",
	230 => X"5451",
	231 => X"509D",
	232 => X"4CCB",
	233 => X"48DD",
	234 => X"44D4",
	235 => X"40B2",
	236 => X"3C78",
	237 => X"3828",
	238 => X"33C3",
	239 => X"2F4C",
	240 => X"2AC3",
	241 => X"262B",
	242 => X"2184",
	243 => X"1CD1",
	244 => X"1814",
	245 => X"134E",
	246 => X"0E80",
	247 => X"09AE",
	others => X"0000"
);

CONSTANT GS3: hex := (
	000 => X"0000",
	001 => X"0527",
	002 => X"0A4C",
	003 => X"0F6D",
	004 => X"1488",
	005 => X"199A",
	006 => X"1EA1",
	007 => X"239C",
	008 => X"2888",
	009 => X"2D63",
	010 => X"322B",
	011 => X"36DE",
	012 => X"3B7B",
	013 => X"3FFF",
	014 => X"4468",
	015 => X"48B5",
	016 => X"4CE4",
	017 => X"50F3",
	018 => X"54E0",
	019 => X"58AA",
	020 => X"5C4F",
	021 => X"5FCE",
	022 => X"6325",
	023 => X"6653",
	024 => X"6956",
	025 => X"6C2E",
	026 => X"6ED9",
	027 => X"7155",
	028 => X"73A3",
	029 => X"75C0",
	030 => X"77AD",
	031 => X"7968",
	032 => X"7AF1",
	033 => X"7C46",
	034 => X"7D68",
	035 => X"7E56",
	036 => X"7F10",
	037 => X"7F94",
	038 => X"7FE4",
	039 => X"7FFF",
	040 => X"7FE4",
	041 => X"7F94",
	042 => X"7F10",
	043 => X"7E56",
	044 => X"7D68",
	045 => X"7C46",
	046 => X"7AF1",
	047 => X"7968",
	048 => X"77AD",
	049 => X"75C0",
	050 => X"73A3",
	051 => X"7155",
	052 => X"6ED9",
	053 => X"6C2E",
	054 => X"6956",
	055 => X"6653",
	056 => X"6325",
	057 => X"5FCE",
	058 => X"5C4F",
	059 => X"58AA",
	060 => X"54E0",
	061 => X"50F3",
	062 => X"4CE4",
	063 => X"48B5",
	064 => X"4468",
	065 => X"3FFF",
	066 => X"3B7B",
	067 => X"36DE",
	068 => X"322B",
	069 => X"2D63",
	070 => X"2888",
	071 => X"239C",
	072 => X"1EA1",
	073 => X"199A",
	074 => X"1488",
	075 => X"0F6D",
	076 => X"0A4C",
	077 => X"0527",
	078 => X"FFFD",
	079 => X"FAD6",
	080 => X"F5B1",
	081 => X"F090",
	082 => X"EB75",
	083 => X"E663",
	084 => X"E15C",
	085 => X"DC61",
	086 => X"D775",
	087 => X"D29A",
	088 => X"CDD2",
	089 => X"C91F",
	090 => X"C482",
	091 => X"BFFE",
	092 => X"BB95",
	093 => X"B748",
	094 => X"B319",
	095 => X"AF0A",
	096 => X"AB1D",
	097 => X"A753",
	098 => X"A3AE",
	099 => X"A02F",
	100 => X"9CD8",
	101 => X"99AA",
	102 => X"96A7",
	103 => X"93CF",
	104 => X"9124",
	105 => X"8EA8",
	106 => X"8C5A",
	107 => X"8A3D",
	108 => X"8850",
	109 => X"8695",
	110 => X"850C",
	111 => X"83B7",
	112 => X"8295",
	113 => X"81A7",
	114 => X"80ED",
	115 => X"8069",
	116 => X"8019",
	117 => X"7FFF",
	118 => X"8019",
	119 => X"8069",
	120 => X"80ED",
	121 => X"81A7",
	122 => X"8295",
	123 => X"83B7",
	124 => X"850C",
	125 => X"8695",
	126 => X"8850",
	127 => X"8A3D",
	128 => X"8C5A",
	129 => X"8EA8",
	130 => X"9124",
	131 => X"93CF",
	132 => X"96A7",
	133 => X"99AA",
	134 => X"9CD8",
	135 => X"A02F",
	136 => X"A3AE",
	137 => X"A753",
	138 => X"AB1D",
	139 => X"AF0A",
	140 => X"B319",
	141 => X"B748",
	142 => X"BB95",
	143 => X"BFFE",
	144 => X"C482",
	145 => X"C91F",
	146 => X"CDD2",
	147 => X"D29A",
	148 => X"D775",
	149 => X"DC61",
	150 => X"E15C",
	151 => X"E663",
	152 => X"EB75",
	153 => X"F090",
	154 => X"F5B1",
	155 => X"FAD6",
	156 => X"0000",
	157 => X"0527",
	158 => X"0A4C",
	159 => X"0F6D",
	160 => X"1488",
	161 => X"199A",
	162 => X"1EA1",
	163 => X"239C",
	164 => X"2888",
	165 => X"2D63",
	166 => X"322B",
	167 => X"36DE",
	168 => X"3B7B",
	169 => X"3FFF",
	170 => X"4468",
	171 => X"48B5",
	172 => X"4CE4",
	173 => X"50F3",
	174 => X"54E0",
	175 => X"58AA",
	176 => X"5C4F",
	177 => X"5FCE",
	178 => X"6325",
	179 => X"6653",
	180 => X"6956",
	181 => X"6C2E",
	182 => X"6ED9",
	183 => X"7155",
	184 => X"73A3",
	185 => X"75C0",
	186 => X"77AD",
	187 => X"7968",
	188 => X"7AF1",
	189 => X"7C46",
	190 => X"7D68",
	191 => X"7E56",
	192 => X"7F10",
	193 => X"7F94",
	194 => X"7FE4",
	195 => X"7FFF",
	196 => X"7FE4",
	197 => X"7F94",
	198 => X"7F10",
	199 => X"7E56",
	200 => X"7D68",
	201 => X"7C46",
	202 => X"7AF1",
	203 => X"7968",
	204 => X"77AD",
	205 => X"75C0",
	206 => X"73A3",
	207 => X"7155",
	208 => X"6ED9",
	209 => X"6C2E",
	210 => X"6956",
	211 => X"6653",
	212 => X"6325",
	213 => X"5FCE",
	214 => X"5C4F",
	215 => X"58AA",
	216 => X"54E0",
	217 => X"50F3",
	218 => X"4CE4",
	219 => X"48B5",
	220 => X"4468",
	221 => X"3FFF",
	222 => X"3B7B",
	223 => X"36DE",
	224 => X"322B",
	225 => X"2D63",
	226 => X"2888",
	227 => X"239C",
	228 => X"1EA1",
	229 => X"199A",
	230 => X"1488",
	231 => X"0F6D",
	232 => X"0A4C",
	233 => X"0527",
	234 => X"FFFD",
	235 => X"FAD6",
	236 => X"F5B1",
	237 => X"F090",
	238 => X"EB75",
	239 => X"E663",
	240 => X"E15C",
	241 => X"DC61",
	242 => X"D775",
	243 => X"D29A",
	244 => X"CDD2",
	245 => X"C91F",
	246 => X"C482",
	247 => X"BFFE",
	others => X"0000"
);

CONSTANT A3: hex := (
	000 => X"0000",
	001 => X"056E",
	002 => X"0ADA",
	003 => X"1041",
	004 => X"15A1",
	005 => X"1AF7",
	006 => X"2040",
	007 => X"257A",
	008 => X"2AA3",
	009 => X"2FB9",
	010 => X"34B8",
	011 => X"399F",
	012 => X"3E6C",
	013 => X"431B",
	014 => X"47AC",
	015 => X"4C1C",
	016 => X"5068",
	017 => X"5490",
	018 => X"5890",
	019 => X"5C68",
	020 => X"6015",
	021 => X"6395",
	022 => X"66E8",
	023 => X"6A0B",
	024 => X"6CFE",
	025 => X"6FBE",
	026 => X"724A",
	027 => X"74A2",
	028 => X"76C4",
	029 => X"78AF",
	030 => X"7A62",
	031 => X"7BDD",
	032 => X"7D1F",
	033 => X"7E27",
	034 => X"7EF5",
	035 => X"7F88",
	036 => X"7FE1",
	037 => X"7FFF",
	038 => X"7FE1",
	039 => X"7F88",
	040 => X"7EF5",
	041 => X"7E27",
	042 => X"7D1F",
	043 => X"7BDD",
	044 => X"7A62",
	045 => X"78AF",
	046 => X"76C4",
	047 => X"74A2",
	048 => X"724A",
	049 => X"6FBE",
	050 => X"6CFE",
	051 => X"6A0B",
	052 => X"66E8",
	053 => X"6395",
	054 => X"6015",
	055 => X"5C68",
	056 => X"5890",
	057 => X"5490",
	058 => X"5068",
	059 => X"4C1C",
	060 => X"47AC",
	061 => X"431B",
	062 => X"3E6C",
	063 => X"399F",
	064 => X"34B8",
	065 => X"2FB9",
	066 => X"2AA3",
	067 => X"257A",
	068 => X"2040",
	069 => X"1AF7",
	070 => X"15A1",
	071 => X"1041",
	072 => X"0ADA",
	073 => X"056E",
	074 => X"0000",
	075 => X"FA8F",
	076 => X"F523",
	077 => X"EFBC",
	078 => X"EA5C",
	079 => X"E506",
	080 => X"DFBD",
	081 => X"DA83",
	082 => X"D55A",
	083 => X"D044",
	084 => X"CB45",
	085 => X"C65E",
	086 => X"C191",
	087 => X"BCE2",
	088 => X"B851",
	089 => X"B3E1",
	090 => X"AF95",
	091 => X"AB6D",
	092 => X"A76D",
	093 => X"A395",
	094 => X"9FE8",
	095 => X"9C68",
	096 => X"9915",
	097 => X"95F2",
	098 => X"92FF",
	099 => X"903F",
	100 => X"8DB3",
	101 => X"8B5B",
	102 => X"8939",
	103 => X"874E",
	104 => X"859B",
	105 => X"8420",
	106 => X"82DE",
	107 => X"81D6",
	108 => X"8108",
	109 => X"8075",
	110 => X"801C",
	111 => X"7FFF",
	112 => X"801C",
	113 => X"8075",
	114 => X"8108",
	115 => X"81D6",
	116 => X"82DE",
	117 => X"8420",
	118 => X"859B",
	119 => X"874E",
	120 => X"8939",
	121 => X"8B5B",
	122 => X"8DB3",
	123 => X"903F",
	124 => X"92FF",
	125 => X"95F2",
	126 => X"9915",
	127 => X"9C68",
	128 => X"9FE8",
	129 => X"A395",
	130 => X"A76D",
	131 => X"AB6D",
	132 => X"AF95",
	133 => X"B3E1",
	134 => X"B851",
	135 => X"BCE2",
	136 => X"C191",
	137 => X"C65E",
	138 => X"CB45",
	139 => X"D044",
	140 => X"D55A",
	141 => X"DA83",
	142 => X"DFBD",
	143 => X"E506",
	144 => X"EA5C",
	145 => X"EFBC",
	146 => X"F523",
	147 => X"FA8F",
	148 => X"0000",
	149 => X"056E",
	150 => X"0ADA",
	151 => X"1041",
	152 => X"15A1",
	153 => X"1AF7",
	154 => X"2040",
	155 => X"257A",
	156 => X"2AA3",
	157 => X"2FB9",
	158 => X"34B8",
	159 => X"399F",
	160 => X"3E6C",
	161 => X"431B",
	162 => X"47AC",
	163 => X"4C1C",
	164 => X"5068",
	165 => X"5490",
	166 => X"5890",
	167 => X"5C68",
	168 => X"6015",
	169 => X"6395",
	170 => X"66E8",
	171 => X"6A0B",
	172 => X"6CFE",
	173 => X"6FBE",
	174 => X"724A",
	175 => X"74A2",
	176 => X"76C4",
	177 => X"78AF",
	178 => X"7A62",
	179 => X"7BDD",
	180 => X"7D1F",
	181 => X"7E27",
	182 => X"7EF5",
	183 => X"7F88",
	184 => X"7FE1",
	185 => X"7FFF",
	186 => X"7FE1",
	187 => X"7F88",
	188 => X"7EF5",
	189 => X"7E27",
	190 => X"7D1F",
	191 => X"7BDD",
	192 => X"7A62",
	193 => X"78AF",
	194 => X"76C4",
	195 => X"74A2",
	196 => X"724A",
	197 => X"6FBE",
	198 => X"6CFE",
	199 => X"6A0B",
	200 => X"66E8",
	201 => X"6395",
	202 => X"6015",
	203 => X"5C68",
	204 => X"5890",
	205 => X"5490",
	206 => X"5068",
	207 => X"4C1C",
	208 => X"47AC",
	209 => X"431B",
	210 => X"3E6C",
	211 => X"399F",
	212 => X"34B8",
	213 => X"2FB9",
	214 => X"2AA3",
	215 => X"257A",
	216 => X"2040",
	217 => X"1AF7",
	218 => X"15A1",
	219 => X"1041",
	220 => X"0ADA",
	221 => X"056E",
	222 => X"FFFD",
	223 => X"FA8F",
	224 => X"F523",
	225 => X"EFBC",
	226 => X"EA5C",
	227 => X"E506",
	228 => X"DFBD",
	229 => X"DA83",
	230 => X"D55A",
	231 => X"D044",
	232 => X"CB45",
	233 => X"C65E",
	234 => X"C191",
	235 => X"BCE2",
	236 => X"B851",
	237 => X"B3E1",
	238 => X"AF95",
	239 => X"AB6D",
	240 => X"A76D",
	241 => X"A395",
	242 => X"9FE8",
	243 => X"9C68",
	244 => X"9915",
	245 => X"95F2",
	246 => X"92FF",
	247 => X"903F",
	others => X"0000"
);

CONSTANT AS3: hex := (
	000 => X"0000",
	001 => X"05C8",
	002 => X"0B8E",
	003 => X"114D",
	004 => X"1704",
	005 => X"1CAE",
	006 => X"224A",
	007 => X"27D3",
	008 => X"2D48",
	009 => X"32A5",
	010 => X"37E8",
	011 => X"3D0D",
	012 => X"4213",
	013 => X"46F5",
	014 => X"4BB3",
	015 => X"5049",
	016 => X"54B5",
	017 => X"58F5",
	018 => X"5D07",
	019 => X"60E7",
	020 => X"6495",
	021 => X"680F",
	022 => X"6B51",
	023 => X"6E5C",
	024 => X"712D",
	025 => X"73C3",
	026 => X"761D",
	027 => X"7838",
	028 => X"7A15",
	029 => X"7BB2",
	030 => X"7D0E",
	031 => X"7E29",
	032 => X"7F02",
	033 => X"7F98",
	034 => X"7FEC",
	035 => X"7FFC",
	036 => X"7FCA",
	037 => X"7F55",
	038 => X"7E9E",
	039 => X"7DA4",
	040 => X"7C68",
	041 => X"7AEC",
	042 => X"792F",
	043 => X"7732",
	044 => X"74F8",
	045 => X"7280",
	046 => X"6FCC",
	047 => X"6CDE",
	048 => X"69B7",
	049 => X"6659",
	050 => X"62C5",
	051 => X"5EFD",
	052 => X"5B04",
	053 => X"56DB",
	054 => X"5285",
	055 => X"4E03",
	056 => X"4959",
	057 => X"4488",
	058 => X"3F94",
	059 => X"3A7E",
	060 => X"354A",
	061 => X"2FFA",
	062 => X"2A91",
	063 => X"2511",
	064 => X"1F7E",
	065 => X"19DB",
	066 => X"142A",
	067 => X"0E6F",
	068 => X"08AC",
	069 => X"02E4",
	070 => X"FD19",
	071 => X"F751",
	072 => X"F18E",
	073 => X"EBD3",
	074 => X"E622",
	075 => X"E07F",
	076 => X"DAEC",
	077 => X"D56C",
	078 => X"D003",
	079 => X"CAB3",
	080 => X"C57F",
	081 => X"C069",
	082 => X"BB75",
	083 => X"B6A4",
	084 => X"B1FA",
	085 => X"AD78",
	086 => X"A922",
	087 => X"A4F9",
	088 => X"A100",
	089 => X"9D38",
	090 => X"99A4",
	091 => X"9646",
	092 => X"931F",
	093 => X"9031",
	094 => X"8D7D",
	095 => X"8B05",
	096 => X"88CB",
	097 => X"86CE",
	098 => X"8511",
	099 => X"8395",
	100 => X"8259",
	101 => X"815F",
	102 => X"80A8",
	103 => X"8033",
	104 => X"8001",
	105 => X"8011",
	106 => X"8065",
	107 => X"80FB",
	108 => X"81D4",
	109 => X"82EF",
	110 => X"844B",
	111 => X"85E8",
	112 => X"87C5",
	113 => X"89E0",
	114 => X"8C3A",
	115 => X"8ED0",
	116 => X"91A1",
	117 => X"94AC",
	118 => X"97EE",
	119 => X"9B68",
	120 => X"9F16",
	121 => X"A2F6",
	122 => X"A708",
	123 => X"AB48",
	124 => X"AFB4",
	125 => X"B44A",
	126 => X"B908",
	127 => X"BDEA",
	128 => X"C2F0",
	129 => X"C815",
	130 => X"CD58",
	131 => X"D2B5",
	132 => X"D82A",
	133 => X"DDB3",
	134 => X"E34F",
	135 => X"E8F9",
	136 => X"EEB0",
	137 => X"F46F",
	138 => X"FA35",
	139 => X"FFFD",
	140 => X"05C8",
	141 => X"0B8E",
	142 => X"114D",
	143 => X"1704",
	144 => X"1CAE",
	145 => X"224A",
	146 => X"27D3",
	147 => X"2D48",
	148 => X"32A5",
	149 => X"37E8",
	150 => X"3D0D",
	151 => X"4213",
	152 => X"46F5",
	153 => X"4BB3",
	154 => X"5049",
	155 => X"54B5",
	156 => X"58F5",
	157 => X"5D07",
	158 => X"60E7",
	159 => X"6495",
	160 => X"680F",
	161 => X"6B51",
	162 => X"6E5C",
	163 => X"712D",
	164 => X"73C3",
	165 => X"761D",
	166 => X"7838",
	167 => X"7A15",
	168 => X"7BB2",
	169 => X"7D0E",
	170 => X"7E29",
	171 => X"7F02",
	172 => X"7F98",
	173 => X"7FEC",
	174 => X"7FFC",
	175 => X"7FCA",
	176 => X"7F55",
	177 => X"7E9E",
	178 => X"7DA4",
	179 => X"7C68",
	180 => X"7AEC",
	181 => X"792F",
	182 => X"7732",
	183 => X"74F8",
	184 => X"7280",
	185 => X"6FCC",
	186 => X"6CDE",
	187 => X"69B7",
	188 => X"6659",
	189 => X"62C5",
	190 => X"5EFD",
	191 => X"5B04",
	192 => X"56DB",
	193 => X"5285",
	194 => X"4E03",
	195 => X"4959",
	196 => X"4488",
	197 => X"3F94",
	198 => X"3A7E",
	199 => X"354A",
	200 => X"2FFA",
	201 => X"2A91",
	202 => X"2511",
	203 => X"1F7E",
	204 => X"19DB",
	205 => X"142A",
	206 => X"0E6F",
	207 => X"08AC",
	208 => X"02E4",
	209 => X"FD19",
	210 => X"F751",
	211 => X"F18E",
	212 => X"EBD3",
	213 => X"E622",
	214 => X"E07F",
	215 => X"DAEC",
	216 => X"D56C",
	217 => X"D003",
	218 => X"CAB3",
	219 => X"C57F",
	220 => X"C069",
	221 => X"BB75",
	222 => X"B6A4",
	223 => X"B1FA",
	224 => X"AD78",
	225 => X"A922",
	226 => X"A4F9",
	227 => X"A100",
	228 => X"9D38",
	229 => X"99A4",
	230 => X"9646",
	231 => X"931F",
	232 => X"9031",
	233 => X"8D7D",
	234 => X"8B05",
	235 => X"88CB",
	236 => X"86CE",
	237 => X"8511",
	238 => X"8395",
	239 => X"8259",
	240 => X"815F",
	241 => X"80A8",
	242 => X"8033",
	243 => X"8001",
	244 => X"8011",
	245 => X"8065",
	246 => X"80FB",
	247 => X"81D4",
	others => X"0000"
);

CONSTANT B3: hex := (
	000 => X"0000",
	001 => X"0623",
	002 => X"0C42",
	003 => X"125A",
	004 => X"1867",
	005 => X"1E66",
	006 => X"2454",
	007 => X"2A2B",
	008 => X"2FEA",
	009 => X"358D",
	010 => X"3B10",
	011 => X"4070",
	012 => X"45AB",
	013 => X"4ABC",
	014 => X"4FA1",
	015 => X"5458",
	016 => X"58DD",
	017 => X"5D2D",
	018 => X"6147",
	019 => X"6527",
	020 => X"68CC",
	021 => X"6C33",
	022 => X"6F5B",
	023 => X"7240",
	024 => X"74E3",
	025 => X"7741",
	026 => X"7958",
	027 => X"7B28",
	028 => X"7CB0",
	029 => X"7DEE",
	030 => X"7EE2",
	031 => X"7F8B",
	032 => X"7FE9",
	033 => X"7FFC",
	034 => X"7FC4",
	035 => X"7F40",
	036 => X"7E71",
	037 => X"7D58",
	038 => X"7BF5",
	039 => X"7A49",
	040 => X"7855",
	041 => X"761B",
	042 => X"739A",
	043 => X"70D6",
	044 => X"6DCF",
	045 => X"6A88",
	046 => X"6701",
	047 => X"633E",
	048 => X"5F41",
	049 => X"5B0C",
	050 => X"56A1",
	051 => X"5203",
	052 => X"4D34",
	053 => X"4839",
	054 => X"4312",
	055 => X"3DC5",
	056 => X"3853",
	057 => X"32BF",
	058 => X"2D0E",
	059 => X"2742",
	060 => X"215F",
	061 => X"1B69",
	062 => X"1562",
	063 => X"0F4F",
	064 => X"0933",
	065 => X"0311",
	066 => X"FCEC",
	067 => X"F6CA",
	068 => X"F0AE",
	069 => X"EA9B",
	070 => X"E494",
	071 => X"DE9E",
	072 => X"D8BB",
	073 => X"D2EF",
	074 => X"CD3E",
	075 => X"C7AA",
	076 => X"C238",
	077 => X"BCEB",
	078 => X"B7C4",
	079 => X"B2C9",
	080 => X"ADFA",
	081 => X"A95C",
	082 => X"A4F1",
	083 => X"A0BC",
	084 => X"9CBF",
	085 => X"98FC",
	086 => X"9575",
	087 => X"922E",
	088 => X"8F27",
	089 => X"8C63",
	090 => X"89E2",
	091 => X"87A8",
	092 => X"85B4",
	093 => X"8408",
	094 => X"82A5",
	095 => X"818C",
	096 => X"80BD",
	097 => X"8039",
	098 => X"8001",
	099 => X"8014",
	100 => X"8072",
	101 => X"811B",
	102 => X"820F",
	103 => X"834D",
	104 => X"84D5",
	105 => X"86A5",
	106 => X"88BC",
	107 => X"8B1A",
	108 => X"8DBD",
	109 => X"90A2",
	110 => X"93CA",
	111 => X"9731",
	112 => X"9AD6",
	113 => X"9EB6",
	114 => X"A2D0",
	115 => X"A720",
	116 => X"ABA5",
	117 => X"B05C",
	118 => X"B541",
	119 => X"BA52",
	120 => X"BF8D",
	121 => X"C4ED",
	122 => X"CA70",
	123 => X"D013",
	124 => X"D5D2",
	125 => X"DBA9",
	126 => X"E197",
	127 => X"E796",
	128 => X"EDA3",
	129 => X"F3BB",
	130 => X"F9DA",
	131 => X"FFFD",
	132 => X"0623",
	133 => X"0C42",
	134 => X"125A",
	135 => X"1867",
	136 => X"1E66",
	137 => X"2454",
	138 => X"2A2B",
	139 => X"2FEA",
	140 => X"358D",
	141 => X"3B10",
	142 => X"4070",
	143 => X"45AB",
	144 => X"4ABC",
	145 => X"4FA1",
	146 => X"5458",
	147 => X"58DD",
	148 => X"5D2D",
	149 => X"6147",
	150 => X"6527",
	151 => X"68CC",
	152 => X"6C33",
	153 => X"6F5B",
	154 => X"7240",
	155 => X"74E3",
	156 => X"7741",
	157 => X"7958",
	158 => X"7B28",
	159 => X"7CB0",
	160 => X"7DEE",
	161 => X"7EE2",
	162 => X"7F8B",
	163 => X"7FE9",
	164 => X"7FFC",
	165 => X"7FC4",
	166 => X"7F40",
	167 => X"7E71",
	168 => X"7D58",
	169 => X"7BF5",
	170 => X"7A49",
	171 => X"7855",
	172 => X"761B",
	173 => X"739A",
	174 => X"70D6",
	175 => X"6DCF",
	176 => X"6A88",
	177 => X"6701",
	178 => X"633E",
	179 => X"5F41",
	180 => X"5B0C",
	181 => X"56A1",
	182 => X"5203",
	183 => X"4D34",
	184 => X"4839",
	185 => X"4312",
	186 => X"3DC5",
	187 => X"3853",
	188 => X"32BF",
	189 => X"2D0E",
	190 => X"2742",
	191 => X"215F",
	192 => X"1B69",
	193 => X"1562",
	194 => X"0F4F",
	195 => X"0933",
	196 => X"0311",
	197 => X"FCEC",
	198 => X"F6CA",
	199 => X"F0AE",
	200 => X"EA9B",
	201 => X"E494",
	202 => X"DE9E",
	203 => X"D8BB",
	204 => X"D2EF",
	205 => X"CD3E",
	206 => X"C7AA",
	207 => X"C238",
	208 => X"BCEB",
	209 => X"B7C4",
	210 => X"B2C9",
	211 => X"ADFA",
	212 => X"A95C",
	213 => X"A4F1",
	214 => X"A0BC",
	215 => X"9CBF",
	216 => X"98FC",
	217 => X"9575",
	218 => X"922E",
	219 => X"8F27",
	220 => X"8C63",
	221 => X"89E2",
	222 => X"87A8",
	223 => X"85B4",
	224 => X"8408",
	225 => X"82A5",
	226 => X"818C",
	227 => X"80BD",
	228 => X"8039",
	229 => X"8001",
	230 => X"8014",
	231 => X"8072",
	232 => X"811B",
	233 => X"820F",
	234 => X"834D",
	235 => X"84D5",
	236 => X"86A5",
	237 => X"88BC",
	238 => X"8B1A",
	239 => X"8DBD",
	240 => X"90A2",
	241 => X"93CA",
	242 => X"9731",
	243 => X"9AD6",
	244 => X"9EB6",
	245 => X"A2D0",
	246 => X"A720",
	247 => X"ABA5",
	others => X"0000"
);

CONSTANT C4: hex := (
	000 => X"0000",
	001 => X"067B",
	002 => X"0CF2",
	003 => X"1361",
	004 => X"19C3",
	005 => X"2015",
	006 => X"2651",
	007 => X"2C74",
	008 => X"3279",
	009 => X"385E",
	010 => X"3E1D",
	011 => X"43B4",
	012 => X"491E",
	013 => X"4E58",
	014 => X"535F",
	015 => X"582F",
	016 => X"5CC5",
	017 => X"611E",
	018 => X"6537",
	019 => X"690D",
	020 => X"6C9F",
	021 => X"6FE9",
	022 => X"72EA",
	023 => X"759F",
	024 => X"7807",
	025 => X"7A20",
	026 => X"7BE8",
	027 => X"7D60",
	028 => X"7E85",
	029 => X"7F56",
	030 => X"7FD4",
	031 => X"7FFF",
	032 => X"7FD4",
	033 => X"7F56",
	034 => X"7E85",
	035 => X"7D60",
	036 => X"7BE8",
	037 => X"7A20",
	038 => X"7807",
	039 => X"759F",
	040 => X"72EA",
	041 => X"6FE9",
	042 => X"6C9F",
	043 => X"690D",
	044 => X"6537",
	045 => X"611E",
	046 => X"5CC5",
	047 => X"582F",
	048 => X"535F",
	049 => X"4E58",
	050 => X"491E",
	051 => X"43B4",
	052 => X"3E1D",
	053 => X"385E",
	054 => X"3279",
	055 => X"2C74",
	056 => X"2651",
	057 => X"2015",
	058 => X"19C3",
	059 => X"1361",
	060 => X"0CF2",
	061 => X"067B",
	062 => X"FFFD",
	063 => X"F982",
	064 => X"F30B",
	065 => X"EC9C",
	066 => X"E63A",
	067 => X"DFE8",
	068 => X"D9AC",
	069 => X"D389",
	070 => X"CD84",
	071 => X"C79F",
	072 => X"C1E0",
	073 => X"BC49",
	074 => X"B6DF",
	075 => X"B1A5",
	076 => X"AC9E",
	077 => X"A7CE",
	078 => X"A338",
	079 => X"9EDF",
	080 => X"9AC6",
	081 => X"96F0",
	082 => X"935E",
	083 => X"9014",
	084 => X"8D13",
	085 => X"8A5E",
	086 => X"87F6",
	087 => X"85DD",
	088 => X"8415",
	089 => X"829D",
	090 => X"8178",
	091 => X"80A7",
	092 => X"8029",
	093 => X"7FFF",
	094 => X"8029",
	095 => X"80A7",
	096 => X"8178",
	097 => X"829D",
	098 => X"8415",
	099 => X"85DD",
	100 => X"87F6",
	101 => X"8A5E",
	102 => X"8D13",
	103 => X"9014",
	104 => X"935E",
	105 => X"96F0",
	106 => X"9AC6",
	107 => X"9EDF",
	108 => X"A338",
	109 => X"A7CE",
	110 => X"AC9E",
	111 => X"B1A5",
	112 => X"B6DF",
	113 => X"BC49",
	114 => X"C1E0",
	115 => X"C79F",
	116 => X"CD84",
	117 => X"D389",
	118 => X"D9AC",
	119 => X"DFE8",
	120 => X"E63A",
	121 => X"EC9C",
	122 => X"F30B",
	123 => X"F982",
	124 => X"FFFD",
	125 => X"067B",
	126 => X"0CF2",
	127 => X"1361",
	128 => X"19C3",
	129 => X"2015",
	130 => X"2651",
	131 => X"2C74",
	132 => X"3279",
	133 => X"385E",
	134 => X"3E1D",
	135 => X"43B4",
	136 => X"491E",
	137 => X"4E58",
	138 => X"535F",
	139 => X"582F",
	140 => X"5CC5",
	141 => X"611E",
	142 => X"6537",
	143 => X"690D",
	144 => X"6C9F",
	145 => X"6FE9",
	146 => X"72EA",
	147 => X"759F",
	148 => X"7807",
	149 => X"7A20",
	150 => X"7BE8",
	151 => X"7D60",
	152 => X"7E85",
	153 => X"7F56",
	154 => X"7FD4",
	155 => X"7FFF",
	156 => X"7FD4",
	157 => X"7F56",
	158 => X"7E85",
	159 => X"7D60",
	160 => X"7BE8",
	161 => X"7A20",
	162 => X"7807",
	163 => X"759F",
	164 => X"72EA",
	165 => X"6FE9",
	166 => X"6C9F",
	167 => X"690D",
	168 => X"6537",
	169 => X"611E",
	170 => X"5CC5",
	171 => X"582F",
	172 => X"535F",
	173 => X"4E58",
	174 => X"491E",
	175 => X"43B4",
	176 => X"3E1D",
	177 => X"385E",
	178 => X"3279",
	179 => X"2C74",
	180 => X"2651",
	181 => X"2015",
	182 => X"19C3",
	183 => X"1361",
	184 => X"0CF2",
	185 => X"067B",
	186 => X"0000",
	187 => X"F982",
	188 => X"F30B",
	189 => X"EC9C",
	190 => X"E63A",
	191 => X"DFE8",
	192 => X"D9AC",
	193 => X"D389",
	194 => X"CD84",
	195 => X"C79F",
	196 => X"C1E0",
	197 => X"BC49",
	198 => X"B6DF",
	199 => X"B1A5",
	200 => X"AC9E",
	201 => X"A7CE",
	202 => X"A338",
	203 => X"9EDF",
	204 => X"9AC6",
	205 => X"96F0",
	206 => X"935E",
	207 => X"9014",
	208 => X"8D13",
	209 => X"8A5E",
	210 => X"87F6",
	211 => X"85DD",
	212 => X"8415",
	213 => X"829D",
	214 => X"8178",
	215 => X"80A7",
	216 => X"8029",
	217 => X"7FFF",
	218 => X"8029",
	219 => X"80A7",
	220 => X"8178",
	221 => X"829D",
	222 => X"8415",
	223 => X"85DD",
	224 => X"87F6",
	225 => X"8A5E",
	226 => X"8D13",
	227 => X"9014",
	228 => X"935E",
	229 => X"96F0",
	230 => X"9AC6",
	231 => X"9EDF",
	232 => X"A338",
	233 => X"A7CE",
	234 => X"AC9E",
	235 => X"B1A5",
	236 => X"B6DF",
	237 => X"BC49",
	238 => X"C1E0",
	239 => X"C79F",
	240 => X"CD84",
	241 => X"D389",
	242 => X"D9AC",
	243 => X"DFE8",
	244 => X"E63A",
	245 => X"EC9C",
	246 => X"F30B",
	247 => X"F982",
	others => X"0000"
);

CONSTANT CS4: hex := (
	000 => X"0000",
	001 => X"06DE",
	002 => X"0DB8",
	003 => X"1488",
	004 => X"1B48",
	005 => X"21F4",
	006 => X"2888",
	007 => X"2EFD",
	008 => X"3550",
	009 => X"3B7B",
	010 => X"417A",
	011 => X"474A",
	012 => X"4CE4",
	013 => X"5246",
	014 => X"576B",
	015 => X"5C4F",
	016 => X"60EF",
	017 => X"6548",
	018 => X"6956",
	019 => X"6D16",
	020 => X"7086",
	021 => X"73A3",
	022 => X"766A",
	023 => X"78DA",
	024 => X"7AF1",
	025 => X"7CAD",
	026 => X"7E0D",
	027 => X"7F10",
	028 => X"7FB5",
	029 => X"7FFC",
	030 => X"7FE4",
	031 => X"7F6E",
	032 => X"7E9A",
	033 => X"7D68",
	034 => X"7BDA",
	035 => X"79F1",
	036 => X"77AD",
	037 => X"7511",
	038 => X"721F",
	039 => X"6ED9",
	040 => X"6B40",
	041 => X"6759",
	042 => X"6325",
	043 => X"5EA8",
	044 => X"59E5",
	045 => X"54E0",
	046 => X"4F9C",
	047 => X"4A1E",
	048 => X"4468",
	049 => X"3E81",
	050 => X"386B",
	051 => X"322B",
	052 => X"2BC6",
	053 => X"2542",
	054 => X"1EA1",
	055 => X"17EA",
	056 => X"1121",
	057 => X"0A4C",
	058 => X"036F",
	059 => X"FC8E",
	060 => X"F5B1",
	061 => X"EEDC",
	062 => X"E813",
	063 => X"E15C",
	064 => X"DABB",
	065 => X"D437",
	066 => X"CDD2",
	067 => X"C792",
	068 => X"C17C",
	069 => X"BB95",
	070 => X"B5DF",
	071 => X"B061",
	072 => X"AB1D",
	073 => X"A618",
	074 => X"A155",
	075 => X"9CD8",
	076 => X"98A4",
	077 => X"94BD",
	078 => X"9124",
	079 => X"8DDE",
	080 => X"8AEC",
	081 => X"8850",
	082 => X"860C",
	083 => X"8423",
	084 => X"8295",
	085 => X"8163",
	086 => X"808F",
	087 => X"8019",
	088 => X"8001",
	089 => X"8048",
	090 => X"80ED",
	091 => X"81F0",
	092 => X"8350",
	093 => X"850C",
	094 => X"8723",
	095 => X"8993",
	096 => X"8C5A",
	097 => X"8F77",
	098 => X"92E7",
	099 => X"96A7",
	100 => X"9AB5",
	101 => X"9F0E",
	102 => X"A3AE",
	103 => X"A892",
	104 => X"ADB7",
	105 => X"B319",
	106 => X"B8B3",
	107 => X"BE83",
	108 => X"C482",
	109 => X"CAAD",
	110 => X"D100",
	111 => X"D775",
	112 => X"DE09",
	113 => X"E4B5",
	114 => X"EB75",
	115 => X"F245",
	116 => X"F91F",
	117 => X"0000",
	118 => X"06DE",
	119 => X"0DB8",
	120 => X"1488",
	121 => X"1B48",
	122 => X"21F4",
	123 => X"2888",
	124 => X"2EFD",
	125 => X"3550",
	126 => X"3B7B",
	127 => X"417A",
	128 => X"474A",
	129 => X"4CE4",
	130 => X"5246",
	131 => X"576B",
	132 => X"5C4F",
	133 => X"60EF",
	134 => X"6548",
	135 => X"6956",
	136 => X"6D16",
	137 => X"7086",
	138 => X"73A3",
	139 => X"766A",
	140 => X"78DA",
	141 => X"7AF1",
	142 => X"7CAD",
	143 => X"7E0D",
	144 => X"7F10",
	145 => X"7FB5",
	146 => X"7FFC",
	147 => X"7FE4",
	148 => X"7F6E",
	149 => X"7E9A",
	150 => X"7D68",
	151 => X"7BDA",
	152 => X"79F1",
	153 => X"77AD",
	154 => X"7511",
	155 => X"721F",
	156 => X"6ED9",
	157 => X"6B40",
	158 => X"6759",
	159 => X"6325",
	160 => X"5EA8",
	161 => X"59E5",
	162 => X"54E0",
	163 => X"4F9C",
	164 => X"4A1E",
	165 => X"4468",
	166 => X"3E81",
	167 => X"386B",
	168 => X"322B",
	169 => X"2BC6",
	170 => X"2542",
	171 => X"1EA1",
	172 => X"17EA",
	173 => X"1121",
	174 => X"0A4C",
	175 => X"036F",
	176 => X"FC8E",
	177 => X"F5B1",
	178 => X"EEDC",
	179 => X"E813",
	180 => X"E15C",
	181 => X"DABB",
	182 => X"D437",
	183 => X"CDD2",
	184 => X"C792",
	185 => X"C17C",
	186 => X"BB95",
	187 => X"B5DF",
	188 => X"B061",
	189 => X"AB1D",
	190 => X"A618",
	191 => X"A155",
	192 => X"9CD8",
	193 => X"98A4",
	194 => X"94BD",
	195 => X"9124",
	196 => X"8DDE",
	197 => X"8AEC",
	198 => X"8850",
	199 => X"860C",
	200 => X"8423",
	201 => X"8295",
	202 => X"8163",
	203 => X"808F",
	204 => X"8019",
	205 => X"8001",
	206 => X"8048",
	207 => X"80ED",
	208 => X"81F0",
	209 => X"8350",
	210 => X"850C",
	211 => X"8723",
	212 => X"8993",
	213 => X"8C5A",
	214 => X"8F77",
	215 => X"92E7",
	216 => X"96A7",
	217 => X"9AB5",
	218 => X"9F0E",
	219 => X"A3AE",
	220 => X"A892",
	221 => X"ADB7",
	222 => X"B319",
	223 => X"B8B3",
	224 => X"BE83",
	225 => X"C482",
	226 => X"CAAD",
	227 => X"D100",
	228 => X"D775",
	229 => X"DE09",
	230 => X"E4B5",
	231 => X"EB75",
	232 => X"F245",
	233 => X"F91F",
	234 => X"0000",
	235 => X"06DE",
	236 => X"0DB8",
	237 => X"1488",
	238 => X"1B48",
	239 => X"21F4",
	240 => X"2888",
	241 => X"2EFD",
	242 => X"3550",
	243 => X"3B7B",
	244 => X"417A",
	245 => X"474A",
	246 => X"4CE4",
	247 => X"5246",
	others => X"0000"
);

CONSTANT D4: hex := (
	000 => X"0000",
	001 => X"074E",
	002 => X"0E97",
	003 => X"15D3",
	004 => X"1CFD",
	005 => X"240F",
	006 => X"2B03",
	007 => X"31D3",
	008 => X"3879",
	009 => X"3EF0",
	010 => X"4533",
	011 => X"4B3B",
	012 => X"5105",
	013 => X"568C",
	014 => X"5BCA",
	015 => X"60BB",
	016 => X"655C",
	017 => X"69A8",
	018 => X"6D9B",
	019 => X"7134",
	020 => X"746D",
	021 => X"7746",
	022 => X"79BB",
	023 => X"7BCA",
	024 => X"7D72",
	025 => X"7EB1",
	026 => X"7F86",
	027 => X"7FF1",
	028 => X"7FF1",
	029 => X"7F86",
	030 => X"7EB1",
	031 => X"7D72",
	032 => X"7BCA",
	033 => X"79BB",
	034 => X"7746",
	035 => X"746D",
	036 => X"7134",
	037 => X"6D9B",
	038 => X"69A8",
	039 => X"655C",
	040 => X"60BB",
	041 => X"5BCA",
	042 => X"568C",
	043 => X"5105",
	044 => X"4B3B",
	045 => X"4533",
	046 => X"3EF0",
	047 => X"3879",
	048 => X"31D3",
	049 => X"2B03",
	050 => X"240F",
	051 => X"1CFD",
	052 => X"15D3",
	053 => X"0E97",
	054 => X"074E",
	055 => X"0000",
	056 => X"F8AF",
	057 => X"F166",
	058 => X"EA2A",
	059 => X"E300",
	060 => X"DBEE",
	061 => X"D4FA",
	062 => X"CE2A",
	063 => X"C784",
	064 => X"C10D",
	065 => X"BACA",
	066 => X"B4C2",
	067 => X"AEF8",
	068 => X"A971",
	069 => X"A433",
	070 => X"9F42",
	071 => X"9AA1",
	072 => X"9655",
	073 => X"9262",
	074 => X"8EC9",
	075 => X"8B90",
	076 => X"88B7",
	077 => X"8642",
	078 => X"8433",
	079 => X"828B",
	080 => X"814C",
	081 => X"8077",
	082 => X"800C",
	083 => X"800C",
	084 => X"8077",
	085 => X"814C",
	086 => X"828B",
	087 => X"8433",
	088 => X"8642",
	089 => X"88B7",
	090 => X"8B90",
	091 => X"8EC9",
	092 => X"9262",
	093 => X"9655",
	094 => X"9AA1",
	095 => X"9F42",
	096 => X"A433",
	097 => X"A971",
	098 => X"AEF8",
	099 => X"B4C2",
	100 => X"BACA",
	101 => X"C10D",
	102 => X"C784",
	103 => X"CE2A",
	104 => X"D4FA",
	105 => X"DBEE",
	106 => X"E300",
	107 => X"EA2A",
	108 => X"F166",
	109 => X"F8AF",
	110 => X"FFFD",
	111 => X"074E",
	112 => X"0E97",
	113 => X"15D3",
	114 => X"1CFD",
	115 => X"240F",
	116 => X"2B03",
	117 => X"31D3",
	118 => X"3879",
	119 => X"3EF0",
	120 => X"4533",
	121 => X"4B3B",
	122 => X"5105",
	123 => X"568C",
	124 => X"5BCA",
	125 => X"60BB",
	126 => X"655C",
	127 => X"69A8",
	128 => X"6D9B",
	129 => X"7134",
	130 => X"746D",
	131 => X"7746",
	132 => X"79BB",
	133 => X"7BCA",
	134 => X"7D72",
	135 => X"7EB1",
	136 => X"7F86",
	137 => X"7FF1",
	138 => X"7FF1",
	139 => X"7F86",
	140 => X"7EB1",
	141 => X"7D72",
	142 => X"7BCA",
	143 => X"79BB",
	144 => X"7746",
	145 => X"746D",
	146 => X"7134",
	147 => X"6D9B",
	148 => X"69A8",
	149 => X"655C",
	150 => X"60BB",
	151 => X"5BCA",
	152 => X"568C",
	153 => X"5105",
	154 => X"4B3B",
	155 => X"4533",
	156 => X"3EF0",
	157 => X"3879",
	158 => X"31D3",
	159 => X"2B03",
	160 => X"240F",
	161 => X"1CFD",
	162 => X"15D3",
	163 => X"0E97",
	164 => X"074E",
	165 => X"0000",
	166 => X"F8AF",
	167 => X"F166",
	168 => X"EA2A",
	169 => X"E300",
	170 => X"DBEE",
	171 => X"D4FA",
	172 => X"CE2A",
	173 => X"C784",
	174 => X"C10D",
	175 => X"BACA",
	176 => X"B4C2",
	177 => X"AEF8",
	178 => X"A971",
	179 => X"A433",
	180 => X"9F42",
	181 => X"9AA1",
	182 => X"9655",
	183 => X"9262",
	184 => X"8EC9",
	185 => X"8B90",
	186 => X"88B7",
	187 => X"8642",
	188 => X"8433",
	189 => X"828B",
	190 => X"814C",
	191 => X"8077",
	192 => X"800C",
	193 => X"800C",
	194 => X"8077",
	195 => X"814C",
	196 => X"828B",
	197 => X"8433",
	198 => X"8642",
	199 => X"88B7",
	200 => X"8B90",
	201 => X"8EC9",
	202 => X"9262",
	203 => X"9655",
	204 => X"9AA1",
	205 => X"9F42",
	206 => X"A433",
	207 => X"A971",
	208 => X"AEF8",
	209 => X"B4C2",
	210 => X"BACA",
	211 => X"C10D",
	212 => X"C784",
	213 => X"CE2A",
	214 => X"D4FA",
	215 => X"DBEE",
	216 => X"E300",
	217 => X"EA2A",
	218 => X"F166",
	219 => X"F8AF",
	220 => X"FFFD",
	221 => X"074E",
	222 => X"0E97",
	223 => X"15D3",
	224 => X"1CFD",
	225 => X"240F",
	226 => X"2B03",
	227 => X"31D3",
	228 => X"3879",
	229 => X"3EF0",
	230 => X"4533",
	231 => X"4B3B",
	232 => X"5105",
	233 => X"568C",
	234 => X"5BCA",
	235 => X"60BB",
	236 => X"655C",
	237 => X"69A8",
	238 => X"6D9B",
	239 => X"7134",
	240 => X"746D",
	241 => X"7746",
	242 => X"79BB",
	243 => X"7BCA",
	244 => X"7D72",
	245 => X"7EB1",
	246 => X"7F86",
	247 => X"7FF1",
	others => X"0000"
);

CONSTANT DS4: hex := (
	000 => X"0000",
	001 => X"07BA",
	002 => X"0F6D",
	003 => X"1712",
	004 => X"1EA1",
	005 => X"2614",
	006 => X"2D63",
	007 => X"3487",
	008 => X"3B7B",
	009 => X"4237",
	010 => X"48B5",
	011 => X"4EF0",
	012 => X"54E0",
	013 => X"5A81",
	014 => X"5FCE",
	015 => X"64C1",
	016 => X"6956",
	017 => X"6D89",
	018 => X"7155",
	019 => X"74B8",
	020 => X"77AD",
	021 => X"7A33",
	022 => X"7C46",
	023 => X"7DE6",
	024 => X"7F10",
	025 => X"7FC3",
	026 => X"7FFF",
	027 => X"7FC3",
	028 => X"7F10",
	029 => X"7DE6",
	030 => X"7C46",
	031 => X"7A33",
	032 => X"77AD",
	033 => X"74B8",
	034 => X"7155",
	035 => X"6D89",
	036 => X"6956",
	037 => X"64C1",
	038 => X"5FCE",
	039 => X"5A81",
	040 => X"54E0",
	041 => X"4EF0",
	042 => X"48B5",
	043 => X"4237",
	044 => X"3B7B",
	045 => X"3487",
	046 => X"2D63",
	047 => X"2614",
	048 => X"1EA1",
	049 => X"1712",
	050 => X"0F6D",
	051 => X"07BA",
	052 => X"0000",
	053 => X"F843",
	054 => X"F090",
	055 => X"E8EB",
	056 => X"E15C",
	057 => X"D9E9",
	058 => X"D29A",
	059 => X"CB76",
	060 => X"C482",
	061 => X"BDC6",
	062 => X"B748",
	063 => X"B10D",
	064 => X"AB1D",
	065 => X"A57C",
	066 => X"A02F",
	067 => X"9B3C",
	068 => X"96A7",
	069 => X"9274",
	070 => X"8EA8",
	071 => X"8B45",
	072 => X"8850",
	073 => X"85CA",
	074 => X"83B7",
	075 => X"8217",
	076 => X"80ED",
	077 => X"803A",
	078 => X"7FFF",
	079 => X"803A",
	080 => X"80ED",
	081 => X"8217",
	082 => X"83B7",
	083 => X"85CA",
	084 => X"8850",
	085 => X"8B45",
	086 => X"8EA8",
	087 => X"9274",
	088 => X"96A7",
	089 => X"9B3C",
	090 => X"A02F",
	091 => X"A57C",
	092 => X"AB1D",
	093 => X"B10D",
	094 => X"B748",
	095 => X"BDC6",
	096 => X"C482",
	097 => X"CB76",
	098 => X"D29A",
	099 => X"D9E9",
	100 => X"E15C",
	101 => X"E8EB",
	102 => X"F090",
	103 => X"F843",
	104 => X"FFFD",
	105 => X"07BA",
	106 => X"0F6D",
	107 => X"1712",
	108 => X"1EA1",
	109 => X"2614",
	110 => X"2D63",
	111 => X"3487",
	112 => X"3B7B",
	113 => X"4237",
	114 => X"48B5",
	115 => X"4EF0",
	116 => X"54E0",
	117 => X"5A81",
	118 => X"5FCE",
	119 => X"64C1",
	120 => X"6956",
	121 => X"6D89",
	122 => X"7155",
	123 => X"74B8",
	124 => X"77AD",
	125 => X"7A33",
	126 => X"7C46",
	127 => X"7DE6",
	128 => X"7F10",
	129 => X"7FC3",
	130 => X"7FFF",
	131 => X"7FC3",
	132 => X"7F10",
	133 => X"7DE6",
	134 => X"7C46",
	135 => X"7A33",
	136 => X"77AD",
	137 => X"74B8",
	138 => X"7155",
	139 => X"6D89",
	140 => X"6956",
	141 => X"64C1",
	142 => X"5FCE",
	143 => X"5A81",
	144 => X"54E0",
	145 => X"4EF0",
	146 => X"48B5",
	147 => X"4237",
	148 => X"3B7B",
	149 => X"3487",
	150 => X"2D63",
	151 => X"2614",
	152 => X"1EA1",
	153 => X"1712",
	154 => X"0F6D",
	155 => X"07BA",
	156 => X"0000",
	157 => X"F843",
	158 => X"F090",
	159 => X"E8EB",
	160 => X"E15C",
	161 => X"D9E9",
	162 => X"D29A",
	163 => X"CB76",
	164 => X"C482",
	165 => X"BDC6",
	166 => X"B748",
	167 => X"B10D",
	168 => X"AB1D",
	169 => X"A57C",
	170 => X"A02F",
	171 => X"9B3C",
	172 => X"96A7",
	173 => X"9274",
	174 => X"8EA8",
	175 => X"8B45",
	176 => X"8850",
	177 => X"85CA",
	178 => X"83B7",
	179 => X"8217",
	180 => X"80ED",
	181 => X"803A",
	182 => X"7FFF",
	183 => X"803A",
	184 => X"80ED",
	185 => X"8217",
	186 => X"83B7",
	187 => X"85CA",
	188 => X"8850",
	189 => X"8B45",
	190 => X"8EA8",
	191 => X"9274",
	192 => X"96A7",
	193 => X"9B3C",
	194 => X"A02F",
	195 => X"A57C",
	196 => X"AB1D",
	197 => X"B10D",
	198 => X"B748",
	199 => X"BDC6",
	200 => X"C482",
	201 => X"CB76",
	202 => X"D29A",
	203 => X"D9E9",
	204 => X"E15C",
	205 => X"E8EB",
	206 => X"F090",
	207 => X"F843",
	208 => X"FFFD",
	209 => X"07BA",
	210 => X"0F6D",
	211 => X"1712",
	212 => X"1EA1",
	213 => X"2614",
	214 => X"2D63",
	215 => X"3487",
	216 => X"3B7B",
	217 => X"4237",
	218 => X"48B5",
	219 => X"4EF0",
	220 => X"54E0",
	221 => X"5A81",
	222 => X"5FCE",
	223 => X"64C1",
	224 => X"6956",
	225 => X"6D89",
	226 => X"7155",
	227 => X"74B8",
	228 => X"77AD",
	229 => X"7A33",
	230 => X"7C46",
	231 => X"7DE6",
	232 => X"7F10",
	233 => X"7FC3",
	234 => X"7FFF",
	235 => X"7FC3",
	236 => X"7F10",
	237 => X"7DE6",
	238 => X"7C46",
	239 => X"7A33",
	240 => X"77AD",
	241 => X"74B8",
	242 => X"7155",
	243 => X"6D89",
	244 => X"6956",
	245 => X"64C1",
	246 => X"5FCE",
	247 => X"5A81",
	others => X"0000"
);

CONSTANT E4: hex := (
	000 => X"0000",
	001 => X"0833",
	002 => X"105E",
	003 => X"1877",
	004 => X"2077",
	005 => X"2855",
	006 => X"3008",
	007 => X"3789",
	008 => X"3ECF",
	009 => X"45D3",
	010 => X"4C8E",
	011 => X"52F8",
	012 => X"590B",
	013 => X"5EC0",
	014 => X"6412",
	015 => X"68FA",
	016 => X"6D74",
	017 => X"717B",
	018 => X"750A",
	019 => X"781E",
	020 => X"7AB4",
	021 => X"7CC9",
	022 => X"7E5A",
	023 => X"7F67",
	024 => X"7FEE",
	025 => X"7FEE",
	026 => X"7F67",
	027 => X"7E5A",
	028 => X"7CC9",
	029 => X"7AB4",
	030 => X"781E",
	031 => X"750A",
	032 => X"717B",
	033 => X"6D74",
	034 => X"68FA",
	035 => X"6412",
	036 => X"5EC0",
	037 => X"590B",
	038 => X"52F8",
	039 => X"4C8E",
	040 => X"45D3",
	041 => X"3ECF",
	042 => X"3789",
	043 => X"3008",
	044 => X"2855",
	045 => X"2077",
	046 => X"1877",
	047 => X"105E",
	048 => X"0833",
	049 => X"0000",
	050 => X"F7CA",
	051 => X"EF9F",
	052 => X"E786",
	053 => X"DF86",
	054 => X"D7A8",
	055 => X"CFF5",
	056 => X"C874",
	057 => X"C12E",
	058 => X"BA2A",
	059 => X"B36F",
	060 => X"AD05",
	061 => X"A6F2",
	062 => X"A13D",
	063 => X"9BEB",
	064 => X"9703",
	065 => X"9289",
	066 => X"8E82",
	067 => X"8AF3",
	068 => X"87DF",
	069 => X"8549",
	070 => X"8334",
	071 => X"81A3",
	072 => X"8096",
	073 => X"800F",
	074 => X"800F",
	075 => X"8096",
	076 => X"81A3",
	077 => X"8334",
	078 => X"8549",
	079 => X"87DF",
	080 => X"8AF3",
	081 => X"8E82",
	082 => X"9289",
	083 => X"9703",
	084 => X"9BEB",
	085 => X"A13D",
	086 => X"A6F2",
	087 => X"AD05",
	088 => X"B36F",
	089 => X"BA2A",
	090 => X"C12E",
	091 => X"C874",
	092 => X"CFF5",
	093 => X"D7A8",
	094 => X"DF86",
	095 => X"E786",
	096 => X"EF9F",
	097 => X"F7CA",
	098 => X"0000",
	099 => X"0833",
	100 => X"105E",
	101 => X"1877",
	102 => X"2077",
	103 => X"2855",
	104 => X"3008",
	105 => X"3789",
	106 => X"3ECF",
	107 => X"45D3",
	108 => X"4C8E",
	109 => X"52F8",
	110 => X"590B",
	111 => X"5EC0",
	112 => X"6412",
	113 => X"68FA",
	114 => X"6D74",
	115 => X"717B",
	116 => X"750A",
	117 => X"781E",
	118 => X"7AB4",
	119 => X"7CC9",
	120 => X"7E5A",
	121 => X"7F67",
	122 => X"7FEE",
	123 => X"7FEE",
	124 => X"7F67",
	125 => X"7E5A",
	126 => X"7CC9",
	127 => X"7AB4",
	128 => X"781E",
	129 => X"750A",
	130 => X"717B",
	131 => X"6D74",
	132 => X"68FA",
	133 => X"6412",
	134 => X"5EC0",
	135 => X"590B",
	136 => X"52F8",
	137 => X"4C8E",
	138 => X"45D3",
	139 => X"3ECF",
	140 => X"3789",
	141 => X"3008",
	142 => X"2855",
	143 => X"2077",
	144 => X"1877",
	145 => X"105E",
	146 => X"0833",
	147 => X"FFFD",
	148 => X"F7CA",
	149 => X"EF9F",
	150 => X"E786",
	151 => X"DF86",
	152 => X"D7A8",
	153 => X"CFF5",
	154 => X"C874",
	155 => X"C12E",
	156 => X"BA2A",
	157 => X"B36F",
	158 => X"AD05",
	159 => X"A6F2",
	160 => X"A13D",
	161 => X"9BEB",
	162 => X"9703",
	163 => X"9289",
	164 => X"8E82",
	165 => X"8AF3",
	166 => X"87DF",
	167 => X"8549",
	168 => X"8334",
	169 => X"81A3",
	170 => X"8096",
	171 => X"800F",
	172 => X"800F",
	173 => X"8096",
	174 => X"81A3",
	175 => X"8334",
	176 => X"8549",
	177 => X"87DF",
	178 => X"8AF3",
	179 => X"8E82",
	180 => X"9289",
	181 => X"9703",
	182 => X"9BEB",
	183 => X"A13D",
	184 => X"A6F2",
	185 => X"AD05",
	186 => X"B36F",
	187 => X"BA2A",
	188 => X"C12E",
	189 => X"C874",
	190 => X"CFF5",
	191 => X"D7A8",
	192 => X"DF86",
	193 => X"E786",
	194 => X"EF9F",
	195 => X"F7CA",
	196 => X"FFFD",
	197 => X"0833",
	198 => X"105E",
	199 => X"1877",
	200 => X"2077",
	201 => X"2855",
	202 => X"3008",
	203 => X"3789",
	204 => X"3ECF",
	205 => X"45D3",
	206 => X"4C8E",
	207 => X"52F8",
	208 => X"590B",
	209 => X"5EC0",
	210 => X"6412",
	211 => X"68FA",
	212 => X"6D74",
	213 => X"717B",
	214 => X"750A",
	215 => X"781E",
	216 => X"7AB4",
	217 => X"7CC9",
	218 => X"7E5A",
	219 => X"7F67",
	220 => X"7FEE",
	221 => X"7FEE",
	222 => X"7F67",
	223 => X"7E5A",
	224 => X"7CC9",
	225 => X"7AB4",
	226 => X"781E",
	227 => X"750A",
	228 => X"717B",
	229 => X"6D74",
	230 => X"68FA",
	231 => X"6412",
	232 => X"5EC0",
	233 => X"590B",
	234 => X"52F8",
	235 => X"4C8E",
	236 => X"45D3",
	237 => X"3ECF",
	238 => X"3789",
	239 => X"3008",
	240 => X"2855",
	241 => X"2077",
	242 => X"1877",
	243 => X"105E",
	244 => X"0833",
	245 => X"0000",
	246 => X"F7CA",
	247 => X"EF9F",
	others => X"0000"
);

CONSTANT F4: hex := (
	000 => X"0000",
	001 => X"08A4",
	002 => X"113E",
	003 => X"19C3",
	004 => X"222B",
	005 => X"2A6B",
	006 => X"3279",
	007 => X"3A4D",
	008 => X"41DC",
	009 => X"491E",
	010 => X"500B",
	011 => X"569B",
	012 => X"5CC5",
	013 => X"6283",
	014 => X"67CD",
	015 => X"6C9F",
	016 => X"70F2",
	017 => X"74C0",
	018 => X"7807",
	019 => X"7AC1",
	020 => X"7CEC",
	021 => X"7E85",
	022 => X"7F8A",
	023 => X"7FFA",
	024 => X"7FD4",
	025 => X"7F1A",
	026 => X"7DCB",
	027 => X"7BE8",
	028 => X"7976",
	029 => X"7675",
	030 => X"72EA",
	031 => X"6ED9",
	032 => X"6A46",
	033 => X"6537",
	034 => X"5FB2",
	035 => X"59BD",
	036 => X"535F",
	037 => X"4CA0",
	038 => X"4587",
	039 => X"3E1D",
	040 => X"366B",
	041 => X"2E79",
	042 => X"2651",
	043 => X"1DFC",
	044 => X"1584",
	045 => X"0CF2",
	046 => X"0452",
	047 => X"FBAB",
	048 => X"F30B",
	049 => X"EA79",
	050 => X"E201",
	051 => X"D9AC",
	052 => X"D184",
	053 => X"C992",
	054 => X"C1E0",
	055 => X"BA76",
	056 => X"B35D",
	057 => X"AC9E",
	058 => X"A640",
	059 => X"A04B",
	060 => X"9AC6",
	061 => X"95B7",
	062 => X"9124",
	063 => X"8D13",
	064 => X"8988",
	065 => X"8687",
	066 => X"8415",
	067 => X"8232",
	068 => X"80E3",
	069 => X"8029",
	070 => X"8003",
	071 => X"8073",
	072 => X"8178",
	073 => X"8311",
	074 => X"853C",
	075 => X"87F6",
	076 => X"8B3D",
	077 => X"8F0B",
	078 => X"935E",
	079 => X"9830",
	080 => X"9D7A",
	081 => X"A338",
	082 => X"A962",
	083 => X"AFF2",
	084 => X"B6DF",
	085 => X"BE21",
	086 => X"C5B0",
	087 => X"CD84",
	088 => X"D592",
	089 => X"DDD2",
	090 => X"E63A",
	091 => X"EEBF",
	092 => X"F759",
	093 => X"0000",
	094 => X"08A4",
	095 => X"113E",
	096 => X"19C3",
	097 => X"222B",
	098 => X"2A6B",
	099 => X"3279",
	100 => X"3A4D",
	101 => X"41DC",
	102 => X"491E",
	103 => X"500B",
	104 => X"569B",
	105 => X"5CC5",
	106 => X"6283",
	107 => X"67CD",
	108 => X"6C9F",
	109 => X"70F2",
	110 => X"74C0",
	111 => X"7807",
	112 => X"7AC1",
	113 => X"7CEC",
	114 => X"7E85",
	115 => X"7F8A",
	116 => X"7FFA",
	117 => X"7FD4",
	118 => X"7F1A",
	119 => X"7DCB",
	120 => X"7BE8",
	121 => X"7976",
	122 => X"7675",
	123 => X"72EA",
	124 => X"6ED9",
	125 => X"6A46",
	126 => X"6537",
	127 => X"5FB2",
	128 => X"59BD",
	129 => X"535F",
	130 => X"4CA0",
	131 => X"4587",
	132 => X"3E1D",
	133 => X"366B",
	134 => X"2E79",
	135 => X"2651",
	136 => X"1DFC",
	137 => X"1584",
	138 => X"0CF2",
	139 => X"0452",
	140 => X"FBAB",
	141 => X"F30B",
	142 => X"EA79",
	143 => X"E201",
	144 => X"D9AC",
	145 => X"D184",
	146 => X"C992",
	147 => X"C1E0",
	148 => X"BA76",
	149 => X"B35D",
	150 => X"AC9E",
	151 => X"A640",
	152 => X"A04B",
	153 => X"9AC6",
	154 => X"95B7",
	155 => X"9124",
	156 => X"8D13",
	157 => X"8988",
	158 => X"8687",
	159 => X"8415",
	160 => X"8232",
	161 => X"80E3",
	162 => X"8029",
	163 => X"8003",
	164 => X"8073",
	165 => X"8178",
	166 => X"8311",
	167 => X"853C",
	168 => X"87F6",
	169 => X"8B3D",
	170 => X"8F0B",
	171 => X"935E",
	172 => X"9830",
	173 => X"9D7A",
	174 => X"A338",
	175 => X"A962",
	176 => X"AFF2",
	177 => X"B6DF",
	178 => X"BE21",
	179 => X"C5B0",
	180 => X"CD84",
	181 => X"D592",
	182 => X"DDD2",
	183 => X"E63A",
	184 => X"EEBF",
	185 => X"F759",
	186 => X"0000",
	187 => X"08A4",
	188 => X"113E",
	189 => X"19C3",
	190 => X"222B",
	191 => X"2A6B",
	192 => X"3279",
	193 => X"3A4D",
	194 => X"41DC",
	195 => X"491E",
	196 => X"500B",
	197 => X"569B",
	198 => X"5CC5",
	199 => X"6283",
	200 => X"67CD",
	201 => X"6C9F",
	202 => X"70F2",
	203 => X"74C0",
	204 => X"7807",
	205 => X"7AC1",
	206 => X"7CEC",
	207 => X"7E85",
	208 => X"7F8A",
	209 => X"7FFA",
	210 => X"7FD4",
	211 => X"7F1A",
	212 => X"7DCB",
	213 => X"7BE8",
	214 => X"7976",
	215 => X"7675",
	216 => X"72EA",
	217 => X"6ED9",
	218 => X"6A46",
	219 => X"6537",
	220 => X"5FB2",
	221 => X"59BD",
	222 => X"535F",
	223 => X"4CA0",
	224 => X"4587",
	225 => X"3E1D",
	226 => X"366B",
	227 => X"2E79",
	228 => X"2651",
	229 => X"1DFC",
	230 => X"1584",
	231 => X"0CF2",
	232 => X"0452",
	233 => X"FBAB",
	234 => X"F30B",
	235 => X"EA79",
	236 => X"E201",
	237 => X"D9AC",
	238 => X"D184",
	239 => X"C992",
	240 => X"C1E0",
	241 => X"BA76",
	242 => X"B35D",
	243 => X"AC9E",
	244 => X"A640",
	245 => X"A04B",
	246 => X"9AC6",
	247 => X"95B7",
	others => X"0000"
);

CONSTANT FS4: hex := (
	000 => X"0000",
	001 => X"0921",
	002 => X"1237",
	003 => X"1B35",
	004 => X"240F",
	005 => X"2CBA",
	006 => X"352B",
	007 => X"3D57",
	008 => X"4533",
	009 => X"4CB4",
	010 => X"53D1",
	011 => X"5A81",
	012 => X"60BB",
	013 => X"6677",
	014 => X"6BAD",
	015 => X"7056",
	016 => X"746D",
	017 => X"77ED",
	018 => X"7ACF",
	019 => X"7D12",
	020 => X"7EB1",
	021 => X"7FAB",
	022 => X"7FFF",
	023 => X"7FAB",
	024 => X"7EB1",
	025 => X"7D12",
	026 => X"7ACF",
	027 => X"77ED",
	028 => X"746D",
	029 => X"7056",
	030 => X"6BAD",
	031 => X"6677",
	032 => X"60BB",
	033 => X"5A81",
	034 => X"53D1",
	035 => X"4CB4",
	036 => X"4533",
	037 => X"3D57",
	038 => X"352B",
	039 => X"2CBA",
	040 => X"240F",
	041 => X"1B35",
	042 => X"1237",
	043 => X"0921",
	044 => X"FFFD",
	045 => X"F6DC",
	046 => X"EDC6",
	047 => X"E4C8",
	048 => X"DBEE",
	049 => X"D343",
	050 => X"CAD2",
	051 => X"C2A6",
	052 => X"BACA",
	053 => X"B349",
	054 => X"AC2C",
	055 => X"A57C",
	056 => X"9F42",
	057 => X"9986",
	058 => X"9450",
	059 => X"8FA7",
	060 => X"8B90",
	061 => X"8810",
	062 => X"852E",
	063 => X"82EB",
	064 => X"814C",
	065 => X"8052",
	066 => X"7FFF",
	067 => X"8052",
	068 => X"814C",
	069 => X"82EB",
	070 => X"852E",
	071 => X"8810",
	072 => X"8B90",
	073 => X"8FA7",
	074 => X"9450",
	075 => X"9986",
	076 => X"9F42",
	077 => X"A57C",
	078 => X"AC2C",
	079 => X"B349",
	080 => X"BACA",
	081 => X"C2A6",
	082 => X"CAD2",
	083 => X"D343",
	084 => X"DBEE",
	085 => X"E4C8",
	086 => X"EDC6",
	087 => X"F6DC",
	088 => X"FFFD",
	089 => X"0921",
	090 => X"1237",
	091 => X"1B35",
	092 => X"240F",
	093 => X"2CBA",
	094 => X"352B",
	095 => X"3D57",
	096 => X"4533",
	097 => X"4CB4",
	098 => X"53D1",
	099 => X"5A81",
	100 => X"60BB",
	101 => X"6677",
	102 => X"6BAD",
	103 => X"7056",
	104 => X"746D",
	105 => X"77ED",
	106 => X"7ACF",
	107 => X"7D12",
	108 => X"7EB1",
	109 => X"7FAB",
	110 => X"7FFF",
	111 => X"7FAB",
	112 => X"7EB1",
	113 => X"7D12",
	114 => X"7ACF",
	115 => X"77ED",
	116 => X"746D",
	117 => X"7056",
	118 => X"6BAD",
	119 => X"6677",
	120 => X"60BB",
	121 => X"5A81",
	122 => X"53D1",
	123 => X"4CB4",
	124 => X"4533",
	125 => X"3D57",
	126 => X"352B",
	127 => X"2CBA",
	128 => X"240F",
	129 => X"1B35",
	130 => X"1237",
	131 => X"0921",
	132 => X"0000",
	133 => X"F6DC",
	134 => X"EDC6",
	135 => X"E4C8",
	136 => X"DBEE",
	137 => X"D343",
	138 => X"CAD2",
	139 => X"C2A6",
	140 => X"BACA",
	141 => X"B349",
	142 => X"AC2C",
	143 => X"A57C",
	144 => X"9F42",
	145 => X"9986",
	146 => X"9450",
	147 => X"8FA7",
	148 => X"8B90",
	149 => X"8810",
	150 => X"852E",
	151 => X"82EB",
	152 => X"814C",
	153 => X"8052",
	154 => X"7FFF",
	155 => X"8052",
	156 => X"814C",
	157 => X"82EB",
	158 => X"852E",
	159 => X"8810",
	160 => X"8B90",
	161 => X"8FA7",
	162 => X"9450",
	163 => X"9986",
	164 => X"9F42",
	165 => X"A57C",
	166 => X"AC2C",
	167 => X"B349",
	168 => X"BACA",
	169 => X"C2A6",
	170 => X"CAD2",
	171 => X"D343",
	172 => X"DBEE",
	173 => X"E4C8",
	174 => X"EDC6",
	175 => X"F6DC",
	176 => X"0000",
	177 => X"0921",
	178 => X"1237",
	179 => X"1B35",
	180 => X"240F",
	181 => X"2CBA",
	182 => X"352B",
	183 => X"3D57",
	184 => X"4533",
	185 => X"4CB4",
	186 => X"53D1",
	187 => X"5A81",
	188 => X"60BB",
	189 => X"6677",
	190 => X"6BAD",
	191 => X"7056",
	192 => X"746D",
	193 => X"77ED",
	194 => X"7ACF",
	195 => X"7D12",
	196 => X"7EB1",
	197 => X"7FAB",
	198 => X"7FFF",
	199 => X"7FAB",
	200 => X"7EB1",
	201 => X"7D12",
	202 => X"7ACF",
	203 => X"77ED",
	204 => X"746D",
	205 => X"7056",
	206 => X"6BAD",
	207 => X"6677",
	208 => X"60BB",
	209 => X"5A81",
	210 => X"53D1",
	211 => X"4CB4",
	212 => X"4533",
	213 => X"3D57",
	214 => X"352B",
	215 => X"2CBA",
	216 => X"240F",
	217 => X"1B35",
	218 => X"1237",
	219 => X"0921",
	220 => X"FFFD",
	221 => X"F6DC",
	222 => X"EDC6",
	223 => X"E4C8",
	224 => X"DBEE",
	225 => X"D343",
	226 => X"CAD2",
	227 => X"C2A6",
	228 => X"BACA",
	229 => X"B349",
	230 => X"AC2C",
	231 => X"A57C",
	232 => X"9F42",
	233 => X"9986",
	234 => X"9450",
	235 => X"8FA7",
	236 => X"8B90",
	237 => X"8810",
	238 => X"852E",
	239 => X"82EB",
	240 => X"814C",
	241 => X"8052",
	242 => X"7FFF",
	243 => X"8052",
	244 => X"814C",
	245 => X"82EB",
	246 => X"852E",
	247 => X"8810",
	others => X"0000"
);

CONSTANT G4: hex := (
	000 => X"0000",
	001 => X"09AE",
	002 => X"134E",
	003 => X"1CD1",
	004 => X"262B",
	005 => X"2F4C",
	006 => X"3828",
	007 => X"40B2",
	008 => X"48DD",
	009 => X"509D",
	010 => X"57E6",
	011 => X"5EAF",
	012 => X"64ED",
	013 => X"6A97",
	014 => X"6FA5",
	015 => X"740F",
	016 => X"77CF",
	017 => X"7ADF",
	018 => X"7D3B",
	019 => X"7EDF",
	020 => X"7FCA",
	021 => X"7FF9",
	022 => X"7F6C",
	023 => X"7E24",
	024 => X"7C24",
	025 => X"796D",
	026 => X"7605",
	027 => X"71EF",
	028 => X"6D32",
	029 => X"67D5",
	030 => X"61E0",
	031 => X"5B5B",
	032 => X"5451",
	033 => X"4CCB",
	034 => X"44D4",
	035 => X"3C78",
	036 => X"33C3",
	037 => X"2AC3",
	038 => X"2184",
	039 => X"1814",
	040 => X"0E80",
	041 => X"04D7",
	042 => X"FB26",
	043 => X"F17D",
	044 => X"E7E9",
	045 => X"DE79",
	046 => X"D53A",
	047 => X"CC3A",
	048 => X"C385",
	049 => X"BB29",
	050 => X"B332",
	051 => X"ABAC",
	052 => X"A4A2",
	053 => X"9E1D",
	054 => X"9828",
	055 => X"92CB",
	056 => X"8E0E",
	057 => X"89F8",
	058 => X"8690",
	059 => X"83D9",
	060 => X"81D9",
	061 => X"8091",
	062 => X"8004",
	063 => X"8033",
	064 => X"811E",
	065 => X"82C2",
	066 => X"851E",
	067 => X"882E",
	068 => X"8BEE",
	069 => X"9058",
	070 => X"9566",
	071 => X"9B10",
	072 => X"A14E",
	073 => X"A817",
	074 => X"AF60",
	075 => X"B720",
	076 => X"BF4B",
	077 => X"C7D5",
	078 => X"D0B1",
	079 => X"D9D2",
	080 => X"E32C",
	081 => X"ECAF",
	082 => X"F64F",
	083 => X"FFFD",
	084 => X"09AE",
	085 => X"134E",
	086 => X"1CD1",
	087 => X"262B",
	088 => X"2F4C",
	089 => X"3828",
	090 => X"40B2",
	091 => X"48DD",
	092 => X"509D",
	093 => X"57E6",
	094 => X"5EAF",
	095 => X"64ED",
	096 => X"6A97",
	097 => X"6FA5",
	098 => X"740F",
	099 => X"77CF",
	100 => X"7ADF",
	101 => X"7D3B",
	102 => X"7EDF",
	103 => X"7FCA",
	104 => X"7FF9",
	105 => X"7F6C",
	106 => X"7E24",
	107 => X"7C24",
	108 => X"796D",
	109 => X"7605",
	110 => X"71EF",
	111 => X"6D32",
	112 => X"67D5",
	113 => X"61E0",
	114 => X"5B5B",
	115 => X"5451",
	116 => X"4CCB",
	117 => X"44D4",
	118 => X"3C78",
	119 => X"33C3",
	120 => X"2AC3",
	121 => X"2184",
	122 => X"1814",
	123 => X"0E80",
	124 => X"04D7",
	125 => X"FB26",
	126 => X"F17D",
	127 => X"E7E9",
	128 => X"DE79",
	129 => X"D53A",
	130 => X"CC3A",
	131 => X"C385",
	132 => X"BB29",
	133 => X"B332",
	134 => X"ABAC",
	135 => X"A4A2",
	136 => X"9E1D",
	137 => X"9828",
	138 => X"92CB",
	139 => X"8E0E",
	140 => X"89F8",
	141 => X"8690",
	142 => X"83D9",
	143 => X"81D9",
	144 => X"8091",
	145 => X"8004",
	146 => X"8033",
	147 => X"811E",
	148 => X"82C2",
	149 => X"851E",
	150 => X"882E",
	151 => X"8BEE",
	152 => X"9058",
	153 => X"9566",
	154 => X"9B10",
	155 => X"A14E",
	156 => X"A817",
	157 => X"AF60",
	158 => X"B720",
	159 => X"BF4B",
	160 => X"C7D5",
	161 => X"D0B1",
	162 => X"D9D2",
	163 => X"E32C",
	164 => X"ECAF",
	165 => X"F64F",
	166 => X"0000",
	167 => X"09AE",
	168 => X"134E",
	169 => X"1CD1",
	170 => X"262B",
	171 => X"2F4C",
	172 => X"3828",
	173 => X"40B2",
	174 => X"48DD",
	175 => X"509D",
	176 => X"57E6",
	177 => X"5EAF",
	178 => X"64ED",
	179 => X"6A97",
	180 => X"6FA5",
	181 => X"740F",
	182 => X"77CF",
	183 => X"7ADF",
	184 => X"7D3B",
	185 => X"7EDF",
	186 => X"7FCA",
	187 => X"7FF9",
	188 => X"7F6C",
	189 => X"7E24",
	190 => X"7C24",
	191 => X"796D",
	192 => X"7605",
	193 => X"71EF",
	194 => X"6D32",
	195 => X"67D5",
	196 => X"61E0",
	197 => X"5B5B",
	198 => X"5451",
	199 => X"4CCB",
	200 => X"44D4",
	201 => X"3C78",
	202 => X"33C3",
	203 => X"2AC3",
	204 => X"2184",
	205 => X"1814",
	206 => X"0E80",
	207 => X"04D7",
	208 => X"FB26",
	209 => X"F17D",
	210 => X"E7E9",
	211 => X"DE79",
	212 => X"D53A",
	213 => X"CC3A",
	214 => X"C385",
	215 => X"BB29",
	216 => X"B332",
	217 => X"ABAC",
	218 => X"A4A2",
	219 => X"9E1D",
	220 => X"9828",
	221 => X"92CB",
	222 => X"8E0E",
	223 => X"89F8",
	224 => X"8690",
	225 => X"83D9",
	226 => X"81D9",
	227 => X"8091",
	228 => X"8004",
	229 => X"8033",
	230 => X"811E",
	231 => X"82C2",
	232 => X"851E",
	233 => X"882E",
	234 => X"8BEE",
	235 => X"9058",
	236 => X"9566",
	237 => X"9B10",
	238 => X"A14E",
	239 => X"A817",
	240 => X"AF60",
	241 => X"B720",
	242 => X"BF4B",
	243 => X"C7D5",
	244 => X"D0B1",
	245 => X"D9D2",
	246 => X"E32C",
	247 => X"ECAF",
	others => X"0000"
);

CONSTANT GS4: hex := (
	000 => X"0000",
	001 => X"0A4C",
	002 => X"1488",
	003 => X"1EA1",
	004 => X"2888",
	005 => X"322B",
	006 => X"3B7B",
	007 => X"4468",
	008 => X"4CE4",
	009 => X"54E0",
	010 => X"5C4F",
	011 => X"6325",
	012 => X"6956",
	013 => X"6ED9",
	014 => X"73A3",
	015 => X"77AD",
	016 => X"7AF1",
	017 => X"7D68",
	018 => X"7F10",
	019 => X"7FE4",
	020 => X"7FE4",
	021 => X"7F10",
	022 => X"7D68",
	023 => X"7AF1",
	024 => X"77AD",
	025 => X"73A3",
	026 => X"6ED9",
	027 => X"6956",
	028 => X"6325",
	029 => X"5C4F",
	030 => X"54E0",
	031 => X"4CE4",
	032 => X"4468",
	033 => X"3B7B",
	034 => X"322B",
	035 => X"2888",
	036 => X"1EA1",
	037 => X"1488",
	038 => X"0A4C",
	039 => X"0000",
	040 => X"F5B1",
	041 => X"EB75",
	042 => X"E15C",
	043 => X"D775",
	044 => X"CDD2",
	045 => X"C482",
	046 => X"BB95",
	047 => X"B319",
	048 => X"AB1D",
	049 => X"A3AE",
	050 => X"9CD8",
	051 => X"96A7",
	052 => X"9124",
	053 => X"8C5A",
	054 => X"8850",
	055 => X"850C",
	056 => X"8295",
	057 => X"80ED",
	058 => X"8019",
	059 => X"8019",
	060 => X"80ED",
	061 => X"8295",
	062 => X"850C",
	063 => X"8850",
	064 => X"8C5A",
	065 => X"9124",
	066 => X"96A7",
	067 => X"9CD8",
	068 => X"A3AE",
	069 => X"AB1D",
	070 => X"B319",
	071 => X"BB95",
	072 => X"C482",
	073 => X"CDD2",
	074 => X"D775",
	075 => X"E15C",
	076 => X"EB75",
	077 => X"F5B1",
	078 => X"0000",
	079 => X"0A4C",
	080 => X"1488",
	081 => X"1EA1",
	082 => X"2888",
	083 => X"322B",
	084 => X"3B7B",
	085 => X"4468",
	086 => X"4CE4",
	087 => X"54E0",
	088 => X"5C4F",
	089 => X"6325",
	090 => X"6956",
	091 => X"6ED9",
	092 => X"73A3",
	093 => X"77AD",
	094 => X"7AF1",
	095 => X"7D68",
	096 => X"7F10",
	097 => X"7FE4",
	098 => X"7FE4",
	099 => X"7F10",
	100 => X"7D68",
	101 => X"7AF1",
	102 => X"77AD",
	103 => X"73A3",
	104 => X"6ED9",
	105 => X"6956",
	106 => X"6325",
	107 => X"5C4F",
	108 => X"54E0",
	109 => X"4CE4",
	110 => X"4468",
	111 => X"3B7B",
	112 => X"322B",
	113 => X"2888",
	114 => X"1EA1",
	115 => X"1488",
	116 => X"0A4C",
	117 => X"FFFD",
	118 => X"F5B1",
	119 => X"EB75",
	120 => X"E15C",
	121 => X"D775",
	122 => X"CDD2",
	123 => X"C482",
	124 => X"BB95",
	125 => X"B319",
	126 => X"AB1D",
	127 => X"A3AE",
	128 => X"9CD8",
	129 => X"96A7",
	130 => X"9124",
	131 => X"8C5A",
	132 => X"8850",
	133 => X"850C",
	134 => X"8295",
	135 => X"80ED",
	136 => X"8019",
	137 => X"8019",
	138 => X"80ED",
	139 => X"8295",
	140 => X"850C",
	141 => X"8850",
	142 => X"8C5A",
	143 => X"9124",
	144 => X"96A7",
	145 => X"9CD8",
	146 => X"A3AE",
	147 => X"AB1D",
	148 => X"B319",
	149 => X"BB95",
	150 => X"C482",
	151 => X"CDD2",
	152 => X"D775",
	153 => X"E15C",
	154 => X"EB75",
	155 => X"F5B1",
	156 => X"0000",
	157 => X"0A4C",
	158 => X"1488",
	159 => X"1EA1",
	160 => X"2888",
	161 => X"322B",
	162 => X"3B7B",
	163 => X"4468",
	164 => X"4CE4",
	165 => X"54E0",
	166 => X"5C4F",
	167 => X"6325",
	168 => X"6956",
	169 => X"6ED9",
	170 => X"73A3",
	171 => X"77AD",
	172 => X"7AF1",
	173 => X"7D68",
	174 => X"7F10",
	175 => X"7FE4",
	176 => X"7FE4",
	177 => X"7F10",
	178 => X"7D68",
	179 => X"7AF1",
	180 => X"77AD",
	181 => X"73A3",
	182 => X"6ED9",
	183 => X"6956",
	184 => X"6325",
	185 => X"5C4F",
	186 => X"54E0",
	187 => X"4CE4",
	188 => X"4468",
	189 => X"3B7B",
	190 => X"322B",
	191 => X"2888",
	192 => X"1EA1",
	193 => X"1488",
	194 => X"0A4C",
	195 => X"FFFD",
	196 => X"F5B1",
	197 => X"EB75",
	198 => X"E15C",
	199 => X"D775",
	200 => X"CDD2",
	201 => X"C482",
	202 => X"BB95",
	203 => X"B319",
	204 => X"AB1D",
	205 => X"A3AE",
	206 => X"9CD8",
	207 => X"96A7",
	208 => X"9124",
	209 => X"8C5A",
	210 => X"8850",
	211 => X"850C",
	212 => X"8295",
	213 => X"80ED",
	214 => X"8019",
	215 => X"8019",
	216 => X"80ED",
	217 => X"8295",
	218 => X"850C",
	219 => X"8850",
	220 => X"8C5A",
	221 => X"9124",
	222 => X"96A7",
	223 => X"9CD8",
	224 => X"A3AE",
	225 => X"AB1D",
	226 => X"B319",
	227 => X"BB95",
	228 => X"C482",
	229 => X"CDD2",
	230 => X"D775",
	231 => X"E15C",
	232 => X"EB75",
	233 => X"F5B1",
	234 => X"0000",
	235 => X"0A4C",
	236 => X"1488",
	237 => X"1EA1",
	238 => X"2888",
	239 => X"322B",
	240 => X"3B7B",
	241 => X"4468",
	242 => X"4CE4",
	243 => X"54E0",
	244 => X"5C4F",
	245 => X"6325",
	246 => X"6956",
	247 => X"6ED9",
	others => X"0000"
);

CONSTANT A4: hex := (
	000 => X"0000",
	001 => X"0ADA",
	002 => X"15A1",
	003 => X"2040",
	004 => X"2AA3",
	005 => X"34B8",
	006 => X"3E6C",
	007 => X"47AC",
	008 => X"5068",
	009 => X"5890",
	010 => X"6015",
	011 => X"66E8",
	012 => X"6CFE",
	013 => X"724A",
	014 => X"76C4",
	015 => X"7A62",
	016 => X"7D1F",
	017 => X"7EF5",
	018 => X"7FE1",
	019 => X"7FE1",
	020 => X"7EF5",
	021 => X"7D1F",
	022 => X"7A62",
	023 => X"76C4",
	024 => X"724A",
	025 => X"6CFE",
	026 => X"66E8",
	027 => X"6015",
	028 => X"5890",
	029 => X"5068",
	030 => X"47AC",
	031 => X"3E6C",
	032 => X"34B8",
	033 => X"2AA3",
	034 => X"2040",
	035 => X"15A1",
	036 => X"0ADA",
	037 => X"FFFD",
	038 => X"F523",
	039 => X"EA5C",
	040 => X"DFBD",
	041 => X"D55A",
	042 => X"CB45",
	043 => X"C191",
	044 => X"B851",
	045 => X"AF95",
	046 => X"A76D",
	047 => X"9FE8",
	048 => X"9915",
	049 => X"92FF",
	050 => X"8DB3",
	051 => X"8939",
	052 => X"859B",
	053 => X"82DE",
	054 => X"8108",
	055 => X"801C",
	056 => X"801C",
	057 => X"8108",
	058 => X"82DE",
	059 => X"859B",
	060 => X"8939",
	061 => X"8DB3",
	062 => X"92FF",
	063 => X"9915",
	064 => X"9FE8",
	065 => X"A76D",
	066 => X"AF95",
	067 => X"B851",
	068 => X"C191",
	069 => X"CB45",
	070 => X"D55A",
	071 => X"DFBD",
	072 => X"EA5C",
	073 => X"F523",
	074 => X"FFFD",
	075 => X"0ADA",
	076 => X"15A1",
	077 => X"2040",
	078 => X"2AA3",
	079 => X"34B8",
	080 => X"3E6C",
	081 => X"47AC",
	082 => X"5068",
	083 => X"5890",
	084 => X"6015",
	085 => X"66E8",
	086 => X"6CFE",
	087 => X"724A",
	088 => X"76C4",
	089 => X"7A62",
	090 => X"7D1F",
	091 => X"7EF5",
	092 => X"7FE1",
	093 => X"7FE1",
	094 => X"7EF5",
	095 => X"7D1F",
	096 => X"7A62",
	097 => X"76C4",
	098 => X"724A",
	099 => X"6CFE",
	100 => X"66E8",
	101 => X"6015",
	102 => X"5890",
	103 => X"5068",
	104 => X"47AC",
	105 => X"3E6C",
	106 => X"34B8",
	107 => X"2AA3",
	108 => X"2040",
	109 => X"15A1",
	110 => X"0ADA",
	111 => X"0000",
	112 => X"F523",
	113 => X"EA5C",
	114 => X"DFBD",
	115 => X"D55A",
	116 => X"CB45",
	117 => X"C191",
	118 => X"B851",
	119 => X"AF95",
	120 => X"A76D",
	121 => X"9FE8",
	122 => X"9915",
	123 => X"92FF",
	124 => X"8DB3",
	125 => X"8939",
	126 => X"859B",
	127 => X"82DE",
	128 => X"8108",
	129 => X"801C",
	130 => X"801C",
	131 => X"8108",
	132 => X"82DE",
	133 => X"859B",
	134 => X"8939",
	135 => X"8DB3",
	136 => X"92FF",
	137 => X"9915",
	138 => X"9FE8",
	139 => X"A76D",
	140 => X"AF95",
	141 => X"B851",
	142 => X"C191",
	143 => X"CB45",
	144 => X"D55A",
	145 => X"DFBD",
	146 => X"EA5C",
	147 => X"F523",
	148 => X"0000",
	149 => X"0ADA",
	150 => X"15A1",
	151 => X"2040",
	152 => X"2AA3",
	153 => X"34B8",
	154 => X"3E6C",
	155 => X"47AC",
	156 => X"5068",
	157 => X"5890",
	158 => X"6015",
	159 => X"66E8",
	160 => X"6CFE",
	161 => X"724A",
	162 => X"76C4",
	163 => X"7A62",
	164 => X"7D1F",
	165 => X"7EF5",
	166 => X"7FE1",
	167 => X"7FE1",
	168 => X"7EF5",
	169 => X"7D1F",
	170 => X"7A62",
	171 => X"76C4",
	172 => X"724A",
	173 => X"6CFE",
	174 => X"66E8",
	175 => X"6015",
	176 => X"5890",
	177 => X"5068",
	178 => X"47AC",
	179 => X"3E6C",
	180 => X"34B8",
	181 => X"2AA3",
	182 => X"2040",
	183 => X"15A1",
	184 => X"0ADA",
	185 => X"FFFD",
	186 => X"F523",
	187 => X"EA5C",
	188 => X"DFBD",
	189 => X"D55A",
	190 => X"CB45",
	191 => X"C191",
	192 => X"B851",
	193 => X"AF95",
	194 => X"A76D",
	195 => X"9FE8",
	196 => X"9915",
	197 => X"92FF",
	198 => X"8DB3",
	199 => X"8939",
	200 => X"859B",
	201 => X"82DE",
	202 => X"8108",
	203 => X"801C",
	204 => X"801C",
	205 => X"8108",
	206 => X"82DE",
	207 => X"859B",
	208 => X"8939",
	209 => X"8DB3",
	210 => X"92FF",
	211 => X"9915",
	212 => X"9FE8",
	213 => X"A76D",
	214 => X"AF95",
	215 => X"B851",
	216 => X"C191",
	217 => X"CB45",
	218 => X"D55A",
	219 => X"DFBD",
	220 => X"EA5C",
	221 => X"F523",
	222 => X"0000",
	223 => X"0ADA",
	224 => X"15A1",
	225 => X"2040",
	226 => X"2AA3",
	227 => X"34B8",
	228 => X"3E6C",
	229 => X"47AC",
	230 => X"5068",
	231 => X"5890",
	232 => X"6015",
	233 => X"66E8",
	234 => X"6CFE",
	235 => X"724A",
	236 => X"76C4",
	237 => X"7A62",
	238 => X"7D1F",
	239 => X"7EF5",
	240 => X"7FE1",
	241 => X"7FE1",
	242 => X"7EF5",
	243 => X"7D1F",
	244 => X"7A62",
	245 => X"76C4",
	246 => X"724A",
	247 => X"6CFE",
	others => X"0000"
);

CONSTANT AS4: hex := (
	000 => X"0000",
	001 => X"0B79",
	002 => X"16DA",
	003 => X"220D",
	004 => X"2CF9",
	005 => X"3789",
	006 => X"41A6",
	007 => X"4B3B",
	008 => X"5436",
	009 => X"5C83",
	010 => X"6412",
	011 => X"6AD2",
	012 => X"70B6",
	013 => X"75B2",
	014 => X"79BB",
	015 => X"7CC9",
	016 => X"7ED6",
	017 => X"7FDE",
	018 => X"7FDE",
	019 => X"7ED6",
	020 => X"7CC9",
	021 => X"79BB",
	022 => X"75B2",
	023 => X"70B6",
	024 => X"6AD2",
	025 => X"6412",
	026 => X"5C83",
	027 => X"5436",
	028 => X"4B3B",
	029 => X"41A6",
	030 => X"3789",
	031 => X"2CF9",
	032 => X"220D",
	033 => X"16DA",
	034 => X"0B79",
	035 => X"0000",
	036 => X"F484",
	037 => X"E923",
	038 => X"DDF0",
	039 => X"D304",
	040 => X"C874",
	041 => X"BE57",
	042 => X"B4C2",
	043 => X"ABC7",
	044 => X"A37A",
	045 => X"9BEB",
	046 => X"952B",
	047 => X"8F47",
	048 => X"8A4B",
	049 => X"8642",
	050 => X"8334",
	051 => X"8127",
	052 => X"801F",
	053 => X"801F",
	054 => X"8127",
	055 => X"8334",
	056 => X"8642",
	057 => X"8A4B",
	058 => X"8F47",
	059 => X"952B",
	060 => X"9BEB",
	061 => X"A37A",
	062 => X"ABC7",
	063 => X"B4C2",
	064 => X"BE57",
	065 => X"C874",
	066 => X"D304",
	067 => X"DDF0",
	068 => X"E923",
	069 => X"F484",
	070 => X"0000",
	071 => X"0B79",
	072 => X"16DA",
	073 => X"220D",
	074 => X"2CF9",
	075 => X"3789",
	076 => X"41A6",
	077 => X"4B3B",
	078 => X"5436",
	079 => X"5C83",
	080 => X"6412",
	081 => X"6AD2",
	082 => X"70B6",
	083 => X"75B2",
	084 => X"79BB",
	085 => X"7CC9",
	086 => X"7ED6",
	087 => X"7FDE",
	088 => X"7FDE",
	089 => X"7ED6",
	090 => X"7CC9",
	091 => X"79BB",
	092 => X"75B2",
	093 => X"70B6",
	094 => X"6AD2",
	095 => X"6412",
	096 => X"5C83",
	097 => X"5436",
	098 => X"4B3B",
	099 => X"41A6",
	100 => X"3789",
	101 => X"2CF9",
	102 => X"220D",
	103 => X"16DA",
	104 => X"0B79",
	105 => X"FFFD",
	106 => X"F484",
	107 => X"E923",
	108 => X"DDF0",
	109 => X"D304",
	110 => X"C874",
	111 => X"BE57",
	112 => X"B4C2",
	113 => X"ABC7",
	114 => X"A37A",
	115 => X"9BEB",
	116 => X"952B",
	117 => X"8F47",
	118 => X"8A4B",
	119 => X"8642",
	120 => X"8334",
	121 => X"8127",
	122 => X"801F",
	123 => X"801F",
	124 => X"8127",
	125 => X"8334",
	126 => X"8642",
	127 => X"8A4B",
	128 => X"8F47",
	129 => X"952B",
	130 => X"9BEB",
	131 => X"A37A",
	132 => X"ABC7",
	133 => X"B4C2",
	134 => X"BE57",
	135 => X"C874",
	136 => X"D304",
	137 => X"DDF0",
	138 => X"E923",
	139 => X"F484",
	140 => X"FFFD",
	141 => X"0B79",
	142 => X"16DA",
	143 => X"220D",
	144 => X"2CF9",
	145 => X"3789",
	146 => X"41A6",
	147 => X"4B3B",
	148 => X"5436",
	149 => X"5C83",
	150 => X"6412",
	151 => X"6AD2",
	152 => X"70B6",
	153 => X"75B2",
	154 => X"79BB",
	155 => X"7CC9",
	156 => X"7ED6",
	157 => X"7FDE",
	158 => X"7FDE",
	159 => X"7ED6",
	160 => X"7CC9",
	161 => X"79BB",
	162 => X"75B2",
	163 => X"70B6",
	164 => X"6AD2",
	165 => X"6412",
	166 => X"5C83",
	167 => X"5436",
	168 => X"4B3B",
	169 => X"41A6",
	170 => X"3789",
	171 => X"2CF9",
	172 => X"220D",
	173 => X"16DA",
	174 => X"0B79",
	175 => X"0000",
	176 => X"F484",
	177 => X"E923",
	178 => X"DDF0",
	179 => X"D304",
	180 => X"C874",
	181 => X"BE57",
	182 => X"B4C2",
	183 => X"ABC7",
	184 => X"A37A",
	185 => X"9BEB",
	186 => X"952B",
	187 => X"8F47",
	188 => X"8A4B",
	189 => X"8642",
	190 => X"8334",
	191 => X"8127",
	192 => X"801F",
	193 => X"801F",
	194 => X"8127",
	195 => X"8334",
	196 => X"8642",
	197 => X"8A4B",
	198 => X"8F47",
	199 => X"952B",
	200 => X"9BEB",
	201 => X"A37A",
	202 => X"ABC7",
	203 => X"B4C2",
	204 => X"BE57",
	205 => X"C874",
	206 => X"D304",
	207 => X"DDF0",
	208 => X"E923",
	209 => X"F484",
	210 => X"FFFD",
	211 => X"0B79",
	212 => X"16DA",
	213 => X"220D",
	214 => X"2CF9",
	215 => X"3789",
	216 => X"41A6",
	217 => X"4B3B",
	218 => X"5436",
	219 => X"5C83",
	220 => X"6412",
	221 => X"6AD2",
	222 => X"70B6",
	223 => X"75B2",
	224 => X"79BB",
	225 => X"7CC9",
	226 => X"7ED6",
	227 => X"7FDE",
	228 => X"7FDE",
	229 => X"7ED6",
	230 => X"7CC9",
	231 => X"79BB",
	232 => X"75B2",
	233 => X"70B6",
	234 => X"6AD2",
	235 => X"6412",
	236 => X"5C83",
	237 => X"5436",
	238 => X"4B3B",
	239 => X"41A6",
	240 => X"3789",
	241 => X"2CF9",
	242 => X"220D",
	243 => X"16DA",
	244 => X"0B79",
	245 => X"0000",
	246 => X"F484",
	247 => X"E923",
	others => X"0000"
);

CONSTANT B4: hex := (
	000 => X"0000",
	001 => X"0C2A",
	002 => X"1839",
	003 => X"240F",
	004 => X"2F92",
	005 => X"3AA6",
	006 => X"4533",
	007 => X"4F1F",
	008 => X"5853",
	009 => X"60BB",
	010 => X"6843",
	011 => X"6ED9",
	012 => X"746D",
	013 => X"78F4",
	014 => X"7C63",
	015 => X"7EB1",
	016 => X"7FD9",
	017 => X"7FD9",
	018 => X"7EB1",
	019 => X"7C63",
	020 => X"78F4",
	021 => X"746D",
	022 => X"6ED9",
	023 => X"6843",
	024 => X"60BB",
	025 => X"5853",
	026 => X"4F1F",
	027 => X"4533",
	028 => X"3AA6",
	029 => X"2F92",
	030 => X"240F",
	031 => X"1839",
	032 => X"0C2A",
	033 => X"FFFD",
	034 => X"F3D3",
	035 => X"E7C4",
	036 => X"DBEE",
	037 => X"D06B",
	038 => X"C557",
	039 => X"BACA",
	040 => X"B0DE",
	041 => X"A7AA",
	042 => X"9F42",
	043 => X"97BA",
	044 => X"9124",
	045 => X"8B90",
	046 => X"8709",
	047 => X"839A",
	048 => X"814C",
	049 => X"8024",
	050 => X"8024",
	051 => X"814C",
	052 => X"839A",
	053 => X"8709",
	054 => X"8B90",
	055 => X"9124",
	056 => X"97BA",
	057 => X"9F42",
	058 => X"A7AA",
	059 => X"B0DE",
	060 => X"BACA",
	061 => X"C557",
	062 => X"D06B",
	063 => X"DBEE",
	064 => X"E7C4",
	065 => X"F3D3",
	066 => X"FFFD",
	067 => X"0C2A",
	068 => X"1839",
	069 => X"240F",
	070 => X"2F92",
	071 => X"3AA6",
	072 => X"4533",
	073 => X"4F1F",
	074 => X"5853",
	075 => X"60BB",
	076 => X"6843",
	077 => X"6ED9",
	078 => X"746D",
	079 => X"78F4",
	080 => X"7C63",
	081 => X"7EB1",
	082 => X"7FD9",
	083 => X"7FD9",
	084 => X"7EB1",
	085 => X"7C63",
	086 => X"78F4",
	087 => X"746D",
	088 => X"6ED9",
	089 => X"6843",
	090 => X"60BB",
	091 => X"5853",
	092 => X"4F1F",
	093 => X"4533",
	094 => X"3AA6",
	095 => X"2F92",
	096 => X"240F",
	097 => X"1839",
	098 => X"0C2A",
	099 => X"0000",
	100 => X"F3D3",
	101 => X"E7C4",
	102 => X"DBEE",
	103 => X"D06B",
	104 => X"C557",
	105 => X"BACA",
	106 => X"B0DE",
	107 => X"A7AA",
	108 => X"9F42",
	109 => X"97BA",
	110 => X"9124",
	111 => X"8B90",
	112 => X"8709",
	113 => X"839A",
	114 => X"814C",
	115 => X"8024",
	116 => X"8024",
	117 => X"814C",
	118 => X"839A",
	119 => X"8709",
	120 => X"8B90",
	121 => X"9124",
	122 => X"97BA",
	123 => X"9F42",
	124 => X"A7AA",
	125 => X"B0DE",
	126 => X"BACA",
	127 => X"C557",
	128 => X"D06B",
	129 => X"DBEE",
	130 => X"E7C4",
	131 => X"F3D3",
	132 => X"0000",
	133 => X"0C2A",
	134 => X"1839",
	135 => X"240F",
	136 => X"2F92",
	137 => X"3AA6",
	138 => X"4533",
	139 => X"4F1F",
	140 => X"5853",
	141 => X"60BB",
	142 => X"6843",
	143 => X"6ED9",
	144 => X"746D",
	145 => X"78F4",
	146 => X"7C63",
	147 => X"7EB1",
	148 => X"7FD9",
	149 => X"7FD9",
	150 => X"7EB1",
	151 => X"7C63",
	152 => X"78F4",
	153 => X"746D",
	154 => X"6ED9",
	155 => X"6843",
	156 => X"60BB",
	157 => X"5853",
	158 => X"4F1F",
	159 => X"4533",
	160 => X"3AA6",
	161 => X"2F92",
	162 => X"240F",
	163 => X"1839",
	164 => X"0C2A",
	165 => X"FFFD",
	166 => X"F3D3",
	167 => X"E7C4",
	168 => X"DBEE",
	169 => X"D06B",
	170 => X"C557",
	171 => X"BACA",
	172 => X"B0DE",
	173 => X"A7AA",
	174 => X"9F42",
	175 => X"97BA",
	176 => X"9124",
	177 => X"8B90",
	178 => X"8709",
	179 => X"839A",
	180 => X"814C",
	181 => X"8024",
	182 => X"8024",
	183 => X"814C",
	184 => X"839A",
	185 => X"8709",
	186 => X"8B90",
	187 => X"9124",
	188 => X"97BA",
	189 => X"9F42",
	190 => X"A7AA",
	191 => X"B0DE",
	192 => X"BACA",
	193 => X"C557",
	194 => X"D06B",
	195 => X"DBEE",
	196 => X"E7C4",
	197 => X"F3D3",
	198 => X"0000",
	199 => X"0C2A",
	200 => X"1839",
	201 => X"240F",
	202 => X"2F92",
	203 => X"3AA6",
	204 => X"4533",
	205 => X"4F1F",
	206 => X"5853",
	207 => X"60BB",
	208 => X"6843",
	209 => X"6ED9",
	210 => X"746D",
	211 => X"78F4",
	212 => X"7C63",
	213 => X"7EB1",
	214 => X"7FD9",
	215 => X"7FD9",
	216 => X"7EB1",
	217 => X"7C63",
	218 => X"78F4",
	219 => X"746D",
	220 => X"6ED9",
	221 => X"6843",
	222 => X"60BB",
	223 => X"5853",
	224 => X"4F1F",
	225 => X"4533",
	226 => X"3AA6",
	227 => X"2F92",
	228 => X"240F",
	229 => X"1839",
	230 => X"0C2A",
	231 => X"FFFD",
	232 => X"F3D3",
	233 => X"E7C4",
	234 => X"DBEE",
	235 => X"D06B",
	236 => X"C557",
	237 => X"BACA",
	238 => X"B0DE",
	239 => X"A7AA",
	240 => X"9F42",
	241 => X"97BA",
	242 => X"9124",
	243 => X"8B90",
	244 => X"8709",
	245 => X"839A",
	246 => X"814C",
	247 => X"8024",
	others => X"0000"
);

CONSTANT C5: hex := (
	000 => X"0000",
	001 => X"0CF2",
	002 => X"19C3",
	003 => X"2651",
	004 => X"3279",
	005 => X"3E1D",
	006 => X"491E",
	007 => X"535F",
	008 => X"5CC5",
	009 => X"6537",
	010 => X"6C9F",
	011 => X"72EA",
	012 => X"7807",
	013 => X"7BE8",
	014 => X"7E85",
	015 => X"7FD4",
	016 => X"7FD4",
	017 => X"7E85",
	018 => X"7BE8",
	019 => X"7807",
	020 => X"72EA",
	021 => X"6C9F",
	022 => X"6537",
	023 => X"5CC5",
	024 => X"535F",
	025 => X"491E",
	026 => X"3E1D",
	027 => X"3279",
	028 => X"2651",
	029 => X"19C3",
	030 => X"0CF2",
	031 => X"FFFD",
	032 => X"F30B",
	033 => X"E63A",
	034 => X"D9AC",
	035 => X"CD84",
	036 => X"C1E0",
	037 => X"B6DF",
	038 => X"AC9E",
	039 => X"A338",
	040 => X"9AC6",
	041 => X"935E",
	042 => X"8D13",
	043 => X"87F6",
	044 => X"8415",
	045 => X"8178",
	046 => X"8029",
	047 => X"8029",
	048 => X"8178",
	049 => X"8415",
	050 => X"87F6",
	051 => X"8D13",
	052 => X"935E",
	053 => X"9AC6",
	054 => X"A338",
	055 => X"AC9E",
	056 => X"B6DF",
	057 => X"C1E0",
	058 => X"CD84",
	059 => X"D9AC",
	060 => X"E63A",
	061 => X"F30B",
	062 => X"0000",
	063 => X"0CF2",
	064 => X"19C3",
	065 => X"2651",
	066 => X"3279",
	067 => X"3E1D",
	068 => X"491E",
	069 => X"535F",
	070 => X"5CC5",
	071 => X"6537",
	072 => X"6C9F",
	073 => X"72EA",
	074 => X"7807",
	075 => X"7BE8",
	076 => X"7E85",
	077 => X"7FD4",
	078 => X"7FD4",
	079 => X"7E85",
	080 => X"7BE8",
	081 => X"7807",
	082 => X"72EA",
	083 => X"6C9F",
	084 => X"6537",
	085 => X"5CC5",
	086 => X"535F",
	087 => X"491E",
	088 => X"3E1D",
	089 => X"3279",
	090 => X"2651",
	091 => X"19C3",
	092 => X"0CF2",
	093 => X"FFFD",
	094 => X"F30B",
	095 => X"E63A",
	096 => X"D9AC",
	097 => X"CD84",
	098 => X"C1E0",
	099 => X"B6DF",
	100 => X"AC9E",
	101 => X"A338",
	102 => X"9AC6",
	103 => X"935E",
	104 => X"8D13",
	105 => X"87F6",
	106 => X"8415",
	107 => X"8178",
	108 => X"8029",
	109 => X"8029",
	110 => X"8178",
	111 => X"8415",
	112 => X"87F6",
	113 => X"8D13",
	114 => X"935E",
	115 => X"9AC6",
	116 => X"A338",
	117 => X"AC9E",
	118 => X"B6DF",
	119 => X"C1E0",
	120 => X"CD84",
	121 => X"D9AC",
	122 => X"E63A",
	123 => X"F30B",
	124 => X"FFFD",
	125 => X"0CF2",
	126 => X"19C3",
	127 => X"2651",
	128 => X"3279",
	129 => X"3E1D",
	130 => X"491E",
	131 => X"535F",
	132 => X"5CC5",
	133 => X"6537",
	134 => X"6C9F",
	135 => X"72EA",
	136 => X"7807",
	137 => X"7BE8",
	138 => X"7E85",
	139 => X"7FD4",
	140 => X"7FD4",
	141 => X"7E85",
	142 => X"7BE8",
	143 => X"7807",
	144 => X"72EA",
	145 => X"6C9F",
	146 => X"6537",
	147 => X"5CC5",
	148 => X"535F",
	149 => X"491E",
	150 => X"3E1D",
	151 => X"3279",
	152 => X"2651",
	153 => X"19C3",
	154 => X"0CF2",
	155 => X"0000",
	156 => X"F30B",
	157 => X"E63A",
	158 => X"D9AC",
	159 => X"CD84",
	160 => X"C1E0",
	161 => X"B6DF",
	162 => X"AC9E",
	163 => X"A338",
	164 => X"9AC6",
	165 => X"935E",
	166 => X"8D13",
	167 => X"87F6",
	168 => X"8415",
	169 => X"8178",
	170 => X"8029",
	171 => X"8029",
	172 => X"8178",
	173 => X"8415",
	174 => X"87F6",
	175 => X"8D13",
	176 => X"935E",
	177 => X"9AC6",
	178 => X"A338",
	179 => X"AC9E",
	180 => X"B6DF",
	181 => X"C1E0",
	182 => X"CD84",
	183 => X"D9AC",
	184 => X"E63A",
	185 => X"F30B",
	186 => X"FFFD",
	187 => X"0CF2",
	188 => X"19C3",
	189 => X"2651",
	190 => X"3279",
	191 => X"3E1D",
	192 => X"491E",
	193 => X"535F",
	194 => X"5CC5",
	195 => X"6537",
	196 => X"6C9F",
	197 => X"72EA",
	198 => X"7807",
	199 => X"7BE8",
	200 => X"7E85",
	201 => X"7FD4",
	202 => X"7FD4",
	203 => X"7E85",
	204 => X"7BE8",
	205 => X"7807",
	206 => X"72EA",
	207 => X"6C9F",
	208 => X"6537",
	209 => X"5CC5",
	210 => X"535F",
	211 => X"491E",
	212 => X"3E1D",
	213 => X"3279",
	214 => X"2651",
	215 => X"19C3",
	216 => X"0CF2",
	217 => X"0000",
	218 => X"F30B",
	219 => X"E63A",
	220 => X"D9AC",
	221 => X"CD84",
	222 => X"C1E0",
	223 => X"B6DF",
	224 => X"AC9E",
	225 => X"A338",
	226 => X"9AC6",
	227 => X"935E",
	228 => X"8D13",
	229 => X"87F6",
	230 => X"8415",
	231 => X"8178",
	232 => X"8029",
	233 => X"8029",
	234 => X"8178",
	235 => X"8415",
	236 => X"87F6",
	237 => X"8D13",
	238 => X"935E",
	239 => X"9AC6",
	240 => X"A338",
	241 => X"AC9E",
	242 => X"B6DF",
	243 => X"C1E0",
	244 => X"CD84",
	245 => X"D9AC",
	246 => X"E63A",
	247 => X"F30B",
	others => X"0000"
);

CONSTANT CS5: hex := (
	000 => X"0000",
	001 => X"0D9A",
	002 => X"1B0E",
	003 => X"2833",
	004 => X"34E3",
	005 => X"40FA",
	006 => X"4C55",
	007 => X"56D2",
	008 => X"6053",
	009 => X"68BD",
	010 => X"6FF7",
	011 => X"75EC",
	012 => X"7A8B",
	013 => X"7DC7",
	014 => X"7F96",
	015 => X"7FF3",
	016 => X"7EDD",
	017 => X"7C56",
	018 => X"7867",
	019 => X"731B",
	020 => X"6C81",
	021 => X"64AC",
	022 => X"5BB4",
	023 => X"51B1",
	024 => X"46C1",
	025 => X"3B04",
	026 => X"2E9C",
	027 => X"21AD",
	028 => X"145C",
	029 => X"06CF",
	030 => X"F92E",
	031 => X"EBA1",
	032 => X"DE50",
	033 => X"D161",
	034 => X"C4F9",
	035 => X"B93C",
	036 => X"AE4C",
	037 => X"A449",
	038 => X"9B51",
	039 => X"937C",
	040 => X"8CE2",
	041 => X"8796",
	042 => X"83A7",
	043 => X"8120",
	044 => X"800A",
	045 => X"8067",
	046 => X"8236",
	047 => X"8572",
	048 => X"8A11",
	049 => X"9006",
	050 => X"9740",
	051 => X"9FAA",
	052 => X"A92B",
	053 => X"B3A8",
	054 => X"BF03",
	055 => X"CB1A",
	056 => X"D7CA",
	057 => X"E4EF",
	058 => X"F263",
	059 => X"0000",
	060 => X"0D9A",
	061 => X"1B0E",
	062 => X"2833",
	063 => X"34E3",
	064 => X"40FA",
	065 => X"4C55",
	066 => X"56D2",
	067 => X"6053",
	068 => X"68BD",
	069 => X"6FF7",
	070 => X"75EC",
	071 => X"7A8B",
	072 => X"7DC7",
	073 => X"7F96",
	074 => X"7FF3",
	075 => X"7EDD",
	076 => X"7C56",
	077 => X"7867",
	078 => X"731B",
	079 => X"6C81",
	080 => X"64AC",
	081 => X"5BB4",
	082 => X"51B1",
	083 => X"46C1",
	084 => X"3B04",
	085 => X"2E9C",
	086 => X"21AD",
	087 => X"145C",
	088 => X"06CF",
	089 => X"F92E",
	090 => X"EBA1",
	091 => X"DE50",
	092 => X"D161",
	093 => X"C4F9",
	094 => X"B93C",
	095 => X"AE4C",
	096 => X"A449",
	097 => X"9B51",
	098 => X"937C",
	099 => X"8CE2",
	100 => X"8796",
	101 => X"83A7",
	102 => X"8120",
	103 => X"800A",
	104 => X"8067",
	105 => X"8236",
	106 => X"8572",
	107 => X"8A11",
	108 => X"9006",
	109 => X"9740",
	110 => X"9FAA",
	111 => X"A92B",
	112 => X"B3A8",
	113 => X"BF03",
	114 => X"CB1A",
	115 => X"D7CA",
	116 => X"E4EF",
	117 => X"F263",
	118 => X"0000",
	119 => X"0D9A",
	120 => X"1B0E",
	121 => X"2833",
	122 => X"34E3",
	123 => X"40FA",
	124 => X"4C55",
	125 => X"56D2",
	126 => X"6053",
	127 => X"68BD",
	128 => X"6FF7",
	129 => X"75EC",
	130 => X"7A8B",
	131 => X"7DC7",
	132 => X"7F96",
	133 => X"7FF3",
	134 => X"7EDD",
	135 => X"7C56",
	136 => X"7867",
	137 => X"731B",
	138 => X"6C81",
	139 => X"64AC",
	140 => X"5BB4",
	141 => X"51B1",
	142 => X"46C1",
	143 => X"3B04",
	144 => X"2E9C",
	145 => X"21AD",
	146 => X"145C",
	147 => X"06CF",
	148 => X"F92E",
	149 => X"EBA1",
	150 => X"DE50",
	151 => X"D161",
	152 => X"C4F9",
	153 => X"B93C",
	154 => X"AE4C",
	155 => X"A449",
	156 => X"9B51",
	157 => X"937C",
	158 => X"8CE2",
	159 => X"8796",
	160 => X"83A7",
	161 => X"8120",
	162 => X"800A",
	163 => X"8067",
	164 => X"8236",
	165 => X"8572",
	166 => X"8A11",
	167 => X"9006",
	168 => X"9740",
	169 => X"9FAA",
	170 => X"A92B",
	171 => X"B3A8",
	172 => X"BF03",
	173 => X"CB1A",
	174 => X"D7CA",
	175 => X"E4EF",
	176 => X"F263",
	177 => X"0000",
	178 => X"0D9A",
	179 => X"1B0E",
	180 => X"2833",
	181 => X"34E3",
	182 => X"40FA",
	183 => X"4C55",
	184 => X"56D2",
	185 => X"6053",
	186 => X"68BD",
	187 => X"6FF7",
	188 => X"75EC",
	189 => X"7A8B",
	190 => X"7DC7",
	191 => X"7F96",
	192 => X"7FF3",
	193 => X"7EDD",
	194 => X"7C56",
	195 => X"7867",
	196 => X"731B",
	197 => X"6C81",
	198 => X"64AC",
	199 => X"5BB4",
	200 => X"51B1",
	201 => X"46C1",
	202 => X"3B04",
	203 => X"2E9C",
	204 => X"21AD",
	205 => X"145C",
	206 => X"06CF",
	207 => X"F92E",
	208 => X"EBA1",
	209 => X"DE50",
	210 => X"D161",
	211 => X"C4F9",
	212 => X"B93C",
	213 => X"AE4C",
	214 => X"A449",
	215 => X"9B51",
	216 => X"937C",
	217 => X"8CE2",
	218 => X"8796",
	219 => X"83A7",
	220 => X"8120",
	221 => X"800A",
	222 => X"8067",
	223 => X"8236",
	224 => X"8572",
	225 => X"8A11",
	226 => X"9006",
	227 => X"9740",
	228 => X"9FAA",
	229 => X"A92B",
	230 => X"B3A8",
	231 => X"BF03",
	232 => X"CB1A",
	233 => X"D7CA",
	234 => X"E4EF",
	235 => X"F263",
	236 => X"0000",
	237 => X"0D9A",
	238 => X"1B0E",
	239 => X"2833",
	240 => X"34E3",
	241 => X"40FA",
	242 => X"4C55",
	243 => X"56D2",
	244 => X"6053",
	245 => X"68BD",
	246 => X"6FF7",
	247 => X"75EC",
	others => X"0000"
);

CONSTANT D5: hex := (
	000 => X"0000",
	001 => X"0E97",
	002 => X"1CFD",
	003 => X"2B03",
	004 => X"3879",
	005 => X"4533",
	006 => X"5105",
	007 => X"5BCA",
	008 => X"655C",
	009 => X"6D9B",
	010 => X"746D",
	011 => X"79BB",
	012 => X"7D72",
	013 => X"7F86",
	014 => X"7FF1",
	015 => X"7EB1",
	016 => X"7BCA",
	017 => X"7746",
	018 => X"7134",
	019 => X"69A8",
	020 => X"60BB",
	021 => X"568C",
	022 => X"4B3B",
	023 => X"3EF0",
	024 => X"31D3",
	025 => X"240F",
	026 => X"15D3",
	027 => X"074E",
	028 => X"F8AF",
	029 => X"EA2A",
	030 => X"DBEE",
	031 => X"CE2A",
	032 => X"C10D",
	033 => X"B4C2",
	034 => X"A971",
	035 => X"9F42",
	036 => X"9655",
	037 => X"8EC9",
	038 => X"88B7",
	039 => X"8433",
	040 => X"814C",
	041 => X"800C",
	042 => X"8077",
	043 => X"828B",
	044 => X"8642",
	045 => X"8B90",
	046 => X"9262",
	047 => X"9AA1",
	048 => X"A433",
	049 => X"AEF8",
	050 => X"BACA",
	051 => X"C784",
	052 => X"D4FA",
	053 => X"E300",
	054 => X"F166",
	055 => X"FFFD",
	056 => X"0E97",
	057 => X"1CFD",
	058 => X"2B03",
	059 => X"3879",
	060 => X"4533",
	061 => X"5105",
	062 => X"5BCA",
	063 => X"655C",
	064 => X"6D9B",
	065 => X"746D",
	066 => X"79BB",
	067 => X"7D72",
	068 => X"7F86",
	069 => X"7FF1",
	070 => X"7EB1",
	071 => X"7BCA",
	072 => X"7746",
	073 => X"7134",
	074 => X"69A8",
	075 => X"60BB",
	076 => X"568C",
	077 => X"4B3B",
	078 => X"3EF0",
	079 => X"31D3",
	080 => X"240F",
	081 => X"15D3",
	082 => X"074E",
	083 => X"F8AF",
	084 => X"EA2A",
	085 => X"DBEE",
	086 => X"CE2A",
	087 => X"C10D",
	088 => X"B4C2",
	089 => X"A971",
	090 => X"9F42",
	091 => X"9655",
	092 => X"8EC9",
	093 => X"88B7",
	094 => X"8433",
	095 => X"814C",
	096 => X"800C",
	097 => X"8077",
	098 => X"828B",
	099 => X"8642",
	100 => X"8B90",
	101 => X"9262",
	102 => X"9AA1",
	103 => X"A433",
	104 => X"AEF8",
	105 => X"BACA",
	106 => X"C784",
	107 => X"D4FA",
	108 => X"E300",
	109 => X"F166",
	110 => X"FFFD",
	111 => X"0E97",
	112 => X"1CFD",
	113 => X"2B03",
	114 => X"3879",
	115 => X"4533",
	116 => X"5105",
	117 => X"5BCA",
	118 => X"655C",
	119 => X"6D9B",
	120 => X"746D",
	121 => X"79BB",
	122 => X"7D72",
	123 => X"7F86",
	124 => X"7FF1",
	125 => X"7EB1",
	126 => X"7BCA",
	127 => X"7746",
	128 => X"7134",
	129 => X"69A8",
	130 => X"60BB",
	131 => X"568C",
	132 => X"4B3B",
	133 => X"3EF0",
	134 => X"31D3",
	135 => X"240F",
	136 => X"15D3",
	137 => X"074E",
	138 => X"F8AF",
	139 => X"EA2A",
	140 => X"DBEE",
	141 => X"CE2A",
	142 => X"C10D",
	143 => X"B4C2",
	144 => X"A971",
	145 => X"9F42",
	146 => X"9655",
	147 => X"8EC9",
	148 => X"88B7",
	149 => X"8433",
	150 => X"814C",
	151 => X"800C",
	152 => X"8077",
	153 => X"828B",
	154 => X"8642",
	155 => X"8B90",
	156 => X"9262",
	157 => X"9AA1",
	158 => X"A433",
	159 => X"AEF8",
	160 => X"BACA",
	161 => X"C784",
	162 => X"D4FA",
	163 => X"E300",
	164 => X"F166",
	165 => X"FFFD",
	166 => X"0E97",
	167 => X"1CFD",
	168 => X"2B03",
	169 => X"3879",
	170 => X"4533",
	171 => X"5105",
	172 => X"5BCA",
	173 => X"655C",
	174 => X"6D9B",
	175 => X"746D",
	176 => X"79BB",
	177 => X"7D72",
	178 => X"7F86",
	179 => X"7FF1",
	180 => X"7EB1",
	181 => X"7BCA",
	182 => X"7746",
	183 => X"7134",
	184 => X"69A8",
	185 => X"60BB",
	186 => X"568C",
	187 => X"4B3B",
	188 => X"3EF0",
	189 => X"31D3",
	190 => X"240F",
	191 => X"15D3",
	192 => X"074E",
	193 => X"F8AF",
	194 => X"EA2A",
	195 => X"DBEE",
	196 => X"CE2A",
	197 => X"C10D",
	198 => X"B4C2",
	199 => X"A971",
	200 => X"9F42",
	201 => X"9655",
	202 => X"8EC9",
	203 => X"88B7",
	204 => X"8433",
	205 => X"814C",
	206 => X"800C",
	207 => X"8077",
	208 => X"828B",
	209 => X"8642",
	210 => X"8B90",
	211 => X"9262",
	212 => X"9AA1",
	213 => X"A433",
	214 => X"AEF8",
	215 => X"BACA",
	216 => X"C784",
	217 => X"D4FA",
	218 => X"E300",
	219 => X"F166",
	220 => X"FFFD",
	221 => X"0E97",
	222 => X"1CFD",
	223 => X"2B03",
	224 => X"3879",
	225 => X"4533",
	226 => X"5105",
	227 => X"5BCA",
	228 => X"655C",
	229 => X"6D9B",
	230 => X"746D",
	231 => X"79BB",
	232 => X"7D72",
	233 => X"7F86",
	234 => X"7FF1",
	235 => X"7EB1",
	236 => X"7BCA",
	237 => X"7746",
	238 => X"7134",
	239 => X"69A8",
	240 => X"60BB",
	241 => X"568C",
	242 => X"4B3B",
	243 => X"3EF0",
	244 => X"31D3",
	245 => X"240F",
	246 => X"15D3",
	247 => X"074E",
	others => X"0000"
);

CONSTANT DS5: hex := (
	000 => X"0000",
	001 => X"0F6D",
	002 => X"1EA1",
	003 => X"2D63",
	004 => X"3B7B",
	005 => X"48B5",
	006 => X"54E0",
	007 => X"5FCE",
	008 => X"6956",
	009 => X"7155",
	010 => X"77AD",
	011 => X"7C46",
	012 => X"7F10",
	013 => X"7FFF",
	014 => X"7F10",
	015 => X"7C46",
	016 => X"77AD",
	017 => X"7155",
	018 => X"6956",
	019 => X"5FCE",
	020 => X"54E0",
	021 => X"48B5",
	022 => X"3B7B",
	023 => X"2D63",
	024 => X"1EA1",
	025 => X"0F6D",
	026 => X"FFFD",
	027 => X"F090",
	028 => X"E15C",
	029 => X"D29A",
	030 => X"C482",
	031 => X"B748",
	032 => X"AB1D",
	033 => X"A02F",
	034 => X"96A7",
	035 => X"8EA8",
	036 => X"8850",
	037 => X"83B7",
	038 => X"80ED",
	039 => X"7FFF",
	040 => X"80ED",
	041 => X"83B7",
	042 => X"8850",
	043 => X"8EA8",
	044 => X"96A7",
	045 => X"A02F",
	046 => X"AB1D",
	047 => X"B748",
	048 => X"C482",
	049 => X"D29A",
	050 => X"E15C",
	051 => X"F090",
	052 => X"FFFD",
	053 => X"0F6D",
	054 => X"1EA1",
	055 => X"2D63",
	056 => X"3B7B",
	057 => X"48B5",
	058 => X"54E0",
	059 => X"5FCE",
	060 => X"6956",
	061 => X"7155",
	062 => X"77AD",
	063 => X"7C46",
	064 => X"7F10",
	065 => X"7FFF",
	066 => X"7F10",
	067 => X"7C46",
	068 => X"77AD",
	069 => X"7155",
	070 => X"6956",
	071 => X"5FCE",
	072 => X"54E0",
	073 => X"48B5",
	074 => X"3B7B",
	075 => X"2D63",
	076 => X"1EA1",
	077 => X"0F6D",
	078 => X"0000",
	079 => X"F090",
	080 => X"E15C",
	081 => X"D29A",
	082 => X"C482",
	083 => X"B748",
	084 => X"AB1D",
	085 => X"A02F",
	086 => X"96A7",
	087 => X"8EA8",
	088 => X"8850",
	089 => X"83B7",
	090 => X"80ED",
	091 => X"7FFF",
	092 => X"80ED",
	093 => X"83B7",
	094 => X"8850",
	095 => X"8EA8",
	096 => X"96A7",
	097 => X"A02F",
	098 => X"AB1D",
	099 => X"B748",
	100 => X"C482",
	101 => X"D29A",
	102 => X"E15C",
	103 => X"F090",
	104 => X"FFFD",
	105 => X"0F6D",
	106 => X"1EA1",
	107 => X"2D63",
	108 => X"3B7B",
	109 => X"48B5",
	110 => X"54E0",
	111 => X"5FCE",
	112 => X"6956",
	113 => X"7155",
	114 => X"77AD",
	115 => X"7C46",
	116 => X"7F10",
	117 => X"7FFF",
	118 => X"7F10",
	119 => X"7C46",
	120 => X"77AD",
	121 => X"7155",
	122 => X"6956",
	123 => X"5FCE",
	124 => X"54E0",
	125 => X"48B5",
	126 => X"3B7B",
	127 => X"2D63",
	128 => X"1EA1",
	129 => X"0F6D",
	130 => X"0000",
	131 => X"F090",
	132 => X"E15C",
	133 => X"D29A",
	134 => X"C482",
	135 => X"B748",
	136 => X"AB1D",
	137 => X"A02F",
	138 => X"96A7",
	139 => X"8EA8",
	140 => X"8850",
	141 => X"83B7",
	142 => X"80ED",
	143 => X"7FFF",
	144 => X"80ED",
	145 => X"83B7",
	146 => X"8850",
	147 => X"8EA8",
	148 => X"96A7",
	149 => X"A02F",
	150 => X"AB1D",
	151 => X"B748",
	152 => X"C482",
	153 => X"D29A",
	154 => X"E15C",
	155 => X"F090",
	156 => X"FFFD",
	157 => X"0F6D",
	158 => X"1EA1",
	159 => X"2D63",
	160 => X"3B7B",
	161 => X"48B5",
	162 => X"54E0",
	163 => X"5FCE",
	164 => X"6956",
	165 => X"7155",
	166 => X"77AD",
	167 => X"7C46",
	168 => X"7F10",
	169 => X"7FFF",
	170 => X"7F10",
	171 => X"7C46",
	172 => X"77AD",
	173 => X"7155",
	174 => X"6956",
	175 => X"5FCE",
	176 => X"54E0",
	177 => X"48B5",
	178 => X"3B7B",
	179 => X"2D63",
	180 => X"1EA1",
	181 => X"0F6D",
	182 => X"0000",
	183 => X"F090",
	184 => X"E15C",
	185 => X"D29A",
	186 => X"C482",
	187 => X"B748",
	188 => X"AB1D",
	189 => X"A02F",
	190 => X"96A7",
	191 => X"8EA8",
	192 => X"8850",
	193 => X"83B7",
	194 => X"80ED",
	195 => X"7FFF",
	196 => X"80ED",
	197 => X"83B7",
	198 => X"8850",
	199 => X"8EA8",
	200 => X"96A7",
	201 => X"A02F",
	202 => X"AB1D",
	203 => X"B748",
	204 => X"C482",
	205 => X"D29A",
	206 => X"E15C",
	207 => X"F090",
	208 => X"FFFD",
	209 => X"0F6D",
	210 => X"1EA1",
	211 => X"2D63",
	212 => X"3B7B",
	213 => X"48B5",
	214 => X"54E0",
	215 => X"5FCE",
	216 => X"6956",
	217 => X"7155",
	218 => X"77AD",
	219 => X"7C46",
	220 => X"7F10",
	221 => X"7FFF",
	222 => X"7F10",
	223 => X"7C46",
	224 => X"77AD",
	225 => X"7155",
	226 => X"6956",
	227 => X"5FCE",
	228 => X"54E0",
	229 => X"48B5",
	230 => X"3B7B",
	231 => X"2D63",
	232 => X"1EA1",
	233 => X"0F6D",
	234 => X"0000",
	235 => X"F090",
	236 => X"E15C",
	237 => X"D29A",
	238 => X"C482",
	239 => X"B748",
	240 => X"AB1D",
	241 => X"A02F",
	242 => X"96A7",
	243 => X"8EA8",
	244 => X"8850",
	245 => X"83B7",
	246 => X"80ED",
	247 => X"7FFF",
	others => X"0000"
);

CONSTANT E5: hex := (
	000 => X"0000",
	001 => X"105E",
	002 => X"2077",
	003 => X"3008",
	004 => X"3ECF",
	005 => X"4C8E",
	006 => X"590B",
	007 => X"6412",
	008 => X"6D74",
	009 => X"750A",
	010 => X"7AB4",
	011 => X"7E5A",
	012 => X"7FEE",
	013 => X"7F67",
	014 => X"7CC9",
	015 => X"781E",
	016 => X"717B",
	017 => X"68FA",
	018 => X"5EC0",
	019 => X"52F8",
	020 => X"45D3",
	021 => X"3789",
	022 => X"2855",
	023 => X"1877",
	024 => X"0833",
	025 => X"F7CA",
	026 => X"E786",
	027 => X"D7A8",
	028 => X"C874",
	029 => X"BA2A",
	030 => X"AD05",
	031 => X"A13D",
	032 => X"9703",
	033 => X"8E82",
	034 => X"87DF",
	035 => X"8334",
	036 => X"8096",
	037 => X"800F",
	038 => X"81A3",
	039 => X"8549",
	040 => X"8AF3",
	041 => X"9289",
	042 => X"9BEB",
	043 => X"A6F2",
	044 => X"B36F",
	045 => X"C12E",
	046 => X"CFF5",
	047 => X"DF86",
	048 => X"EF9F",
	049 => X"FFFD",
	050 => X"105E",
	051 => X"2077",
	052 => X"3008",
	053 => X"3ECF",
	054 => X"4C8E",
	055 => X"590B",
	056 => X"6412",
	057 => X"6D74",
	058 => X"750A",
	059 => X"7AB4",
	060 => X"7E5A",
	061 => X"7FEE",
	062 => X"7F67",
	063 => X"7CC9",
	064 => X"781E",
	065 => X"717B",
	066 => X"68FA",
	067 => X"5EC0",
	068 => X"52F8",
	069 => X"45D3",
	070 => X"3789",
	071 => X"2855",
	072 => X"1877",
	073 => X"0833",
	074 => X"F7CA",
	075 => X"E786",
	076 => X"D7A8",
	077 => X"C874",
	078 => X"BA2A",
	079 => X"AD05",
	080 => X"A13D",
	081 => X"9703",
	082 => X"8E82",
	083 => X"87DF",
	084 => X"8334",
	085 => X"8096",
	086 => X"800F",
	087 => X"81A3",
	088 => X"8549",
	089 => X"8AF3",
	090 => X"9289",
	091 => X"9BEB",
	092 => X"A6F2",
	093 => X"B36F",
	094 => X"C12E",
	095 => X"CFF5",
	096 => X"DF86",
	097 => X"EF9F",
	098 => X"0000",
	099 => X"105E",
	100 => X"2077",
	101 => X"3008",
	102 => X"3ECF",
	103 => X"4C8E",
	104 => X"590B",
	105 => X"6412",
	106 => X"6D74",
	107 => X"750A",
	108 => X"7AB4",
	109 => X"7E5A",
	110 => X"7FEE",
	111 => X"7F67",
	112 => X"7CC9",
	113 => X"781E",
	114 => X"717B",
	115 => X"68FA",
	116 => X"5EC0",
	117 => X"52F8",
	118 => X"45D3",
	119 => X"3789",
	120 => X"2855",
	121 => X"1877",
	122 => X"0833",
	123 => X"F7CA",
	124 => X"E786",
	125 => X"D7A8",
	126 => X"C874",
	127 => X"BA2A",
	128 => X"AD05",
	129 => X"A13D",
	130 => X"9703",
	131 => X"8E82",
	132 => X"87DF",
	133 => X"8334",
	134 => X"8096",
	135 => X"800F",
	136 => X"81A3",
	137 => X"8549",
	138 => X"8AF3",
	139 => X"9289",
	140 => X"9BEB",
	141 => X"A6F2",
	142 => X"B36F",
	143 => X"C12E",
	144 => X"CFF5",
	145 => X"DF86",
	146 => X"EF9F",
	147 => X"0000",
	148 => X"105E",
	149 => X"2077",
	150 => X"3008",
	151 => X"3ECF",
	152 => X"4C8E",
	153 => X"590B",
	154 => X"6412",
	155 => X"6D74",
	156 => X"750A",
	157 => X"7AB4",
	158 => X"7E5A",
	159 => X"7FEE",
	160 => X"7F67",
	161 => X"7CC9",
	162 => X"781E",
	163 => X"717B",
	164 => X"68FA",
	165 => X"5EC0",
	166 => X"52F8",
	167 => X"45D3",
	168 => X"3789",
	169 => X"2855",
	170 => X"1877",
	171 => X"0833",
	172 => X"F7CA",
	173 => X"E786",
	174 => X"D7A8",
	175 => X"C874",
	176 => X"BA2A",
	177 => X"AD05",
	178 => X"A13D",
	179 => X"9703",
	180 => X"8E82",
	181 => X"87DF",
	182 => X"8334",
	183 => X"8096",
	184 => X"800F",
	185 => X"81A3",
	186 => X"8549",
	187 => X"8AF3",
	188 => X"9289",
	189 => X"9BEB",
	190 => X"A6F2",
	191 => X"B36F",
	192 => X"C12E",
	193 => X"CFF5",
	194 => X"DF86",
	195 => X"EF9F",
	196 => X"FFFD",
	197 => X"105E",
	198 => X"2077",
	199 => X"3008",
	200 => X"3ECF",
	201 => X"4C8E",
	202 => X"590B",
	203 => X"6412",
	204 => X"6D74",
	205 => X"750A",
	206 => X"7AB4",
	207 => X"7E5A",
	208 => X"7FEE",
	209 => X"7F67",
	210 => X"7CC9",
	211 => X"781E",
	212 => X"717B",
	213 => X"68FA",
	214 => X"5EC0",
	215 => X"52F8",
	216 => X"45D3",
	217 => X"3789",
	218 => X"2855",
	219 => X"1877",
	220 => X"0833",
	221 => X"F7CA",
	222 => X"E786",
	223 => X"D7A8",
	224 => X"C874",
	225 => X"BA2A",
	226 => X"AD05",
	227 => X"A13D",
	228 => X"9703",
	229 => X"8E82",
	230 => X"87DF",
	231 => X"8334",
	232 => X"8096",
	233 => X"800F",
	234 => X"81A3",
	235 => X"8549",
	236 => X"8AF3",
	237 => X"9289",
	238 => X"9BEB",
	239 => X"A6F2",
	240 => X"B36F",
	241 => X"C12E",
	242 => X"CFF5",
	243 => X"DF86",
	244 => X"EF9F",
	245 => X"FFFD",
	246 => X"105E",
	247 => X"2077",
	others => X"0000"
);

CONSTANT F5: hex := (
	000 => X"0000",
	001 => X"110F",
	002 => X"21D0",
	003 => X"31F7",
	004 => X"413A",
	005 => X"4F53",
	006 => X"5C01",
	007 => X"670B",
	008 => X"703F",
	009 => X"7771",
	010 => X"7C82",
	011 => X"7F5A",
	012 => X"7FEC",
	013 => X"7E36",
	014 => X"7A3F",
	015 => X"741A",
	016 => X"6BE3",
	017 => X"61BE",
	018 => X"55DB",
	019 => X"4870",
	020 => X"39BA",
	021 => X"29FC",
	022 => X"197E",
	023 => X"088C",
	024 => X"F771",
	025 => X"E67F",
	026 => X"D601",
	027 => X"C643",
	028 => X"B78D",
	029 => X"AA22",
	030 => X"9E3F",
	031 => X"941A",
	032 => X"8BE3",
	033 => X"85BE",
	034 => X"81C7",
	035 => X"8011",
	036 => X"80A3",
	037 => X"837B",
	038 => X"888C",
	039 => X"8FBE",
	040 => X"98F2",
	041 => X"A3FC",
	042 => X"B0AA",
	043 => X"BEC3",
	044 => X"CE06",
	045 => X"DE2D",
	046 => X"EEEE",
	047 => X"0000",
	048 => X"110F",
	049 => X"21D0",
	050 => X"31F7",
	051 => X"413A",
	052 => X"4F53",
	053 => X"5C01",
	054 => X"670B",
	055 => X"703F",
	056 => X"7771",
	057 => X"7C82",
	058 => X"7F5A",
	059 => X"7FEC",
	060 => X"7E36",
	061 => X"7A3F",
	062 => X"741A",
	063 => X"6BE3",
	064 => X"61BE",
	065 => X"55DB",
	066 => X"4870",
	067 => X"39BA",
	068 => X"29FC",
	069 => X"197E",
	070 => X"088C",
	071 => X"F771",
	072 => X"E67F",
	073 => X"D601",
	074 => X"C643",
	075 => X"B78D",
	076 => X"AA22",
	077 => X"9E3F",
	078 => X"941A",
	079 => X"8BE3",
	080 => X"85BE",
	081 => X"81C7",
	082 => X"8011",
	083 => X"80A3",
	084 => X"837B",
	085 => X"888C",
	086 => X"8FBE",
	087 => X"98F2",
	088 => X"A3FC",
	089 => X"B0AA",
	090 => X"BEC3",
	091 => X"CE06",
	092 => X"DE2D",
	093 => X"EEEE",
	094 => X"0000",
	095 => X"110F",
	096 => X"21D0",
	097 => X"31F7",
	098 => X"413A",
	099 => X"4F53",
	100 => X"5C01",
	101 => X"670B",
	102 => X"703F",
	103 => X"7771",
	104 => X"7C82",
	105 => X"7F5A",
	106 => X"7FEC",
	107 => X"7E36",
	108 => X"7A3F",
	109 => X"741A",
	110 => X"6BE3",
	111 => X"61BE",
	112 => X"55DB",
	113 => X"4870",
	114 => X"39BA",
	115 => X"29FC",
	116 => X"197E",
	117 => X"088C",
	118 => X"F771",
	119 => X"E67F",
	120 => X"D601",
	121 => X"C643",
	122 => X"B78D",
	123 => X"AA22",
	124 => X"9E3F",
	125 => X"941A",
	126 => X"8BE3",
	127 => X"85BE",
	128 => X"81C7",
	129 => X"8011",
	130 => X"80A3",
	131 => X"837B",
	132 => X"888C",
	133 => X"8FBE",
	134 => X"98F2",
	135 => X"A3FC",
	136 => X"B0AA",
	137 => X"BEC3",
	138 => X"CE06",
	139 => X"DE2D",
	140 => X"EEEE",
	141 => X"0000",
	142 => X"110F",
	143 => X"21D0",
	144 => X"31F7",
	145 => X"413A",
	146 => X"4F53",
	147 => X"5C01",
	148 => X"670B",
	149 => X"703F",
	150 => X"7771",
	151 => X"7C82",
	152 => X"7F5A",
	153 => X"7FEC",
	154 => X"7E36",
	155 => X"7A3F",
	156 => X"741A",
	157 => X"6BE3",
	158 => X"61BE",
	159 => X"55DB",
	160 => X"4870",
	161 => X"39BA",
	162 => X"29FC",
	163 => X"197E",
	164 => X"088C",
	165 => X"F771",
	166 => X"E67F",
	167 => X"D601",
	168 => X"C643",
	169 => X"B78D",
	170 => X"AA22",
	171 => X"9E3F",
	172 => X"941A",
	173 => X"8BE3",
	174 => X"85BE",
	175 => X"81C7",
	176 => X"8011",
	177 => X"80A3",
	178 => X"837B",
	179 => X"888C",
	180 => X"8FBE",
	181 => X"98F2",
	182 => X"A3FC",
	183 => X"B0AA",
	184 => X"BEC3",
	185 => X"CE06",
	186 => X"DE2D",
	187 => X"EEEE",
	188 => X"0000",
	189 => X"110F",
	190 => X"21D0",
	191 => X"31F7",
	192 => X"413A",
	193 => X"4F53",
	194 => X"5C01",
	195 => X"670B",
	196 => X"703F",
	197 => X"7771",
	198 => X"7C82",
	199 => X"7F5A",
	200 => X"7FEC",
	201 => X"7E36",
	202 => X"7A3F",
	203 => X"741A",
	204 => X"6BE3",
	205 => X"61BE",
	206 => X"55DB",
	207 => X"4870",
	208 => X"39BA",
	209 => X"29FC",
	210 => X"197E",
	211 => X"088C",
	212 => X"F771",
	213 => X"E67F",
	214 => X"D601",
	215 => X"C643",
	216 => X"B78D",
	217 => X"AA22",
	218 => X"9E3F",
	219 => X"941A",
	220 => X"8BE3",
	221 => X"85BE",
	222 => X"81C7",
	223 => X"8011",
	224 => X"80A3",
	225 => X"837B",
	226 => X"888C",
	227 => X"8FBE",
	228 => X"98F2",
	229 => X"A3FC",
	230 => X"B0AA",
	231 => X"BEC3",
	232 => X"CE06",
	233 => X"DE2D",
	234 => X"EEEE",
	235 => X"0000",
	236 => X"110F",
	237 => X"21D0",
	238 => X"31F7",
	239 => X"413A",
	240 => X"4F53",
	241 => X"5C01",
	242 => X"670B",
	243 => X"703F",
	244 => X"7771",
	245 => X"7C82",
	246 => X"7F5A",
	247 => X"7FEC",
	others => X"0000"
);

CONSTANT FS5: hex := (
	000 => X"0000",
	001 => X"1237",
	002 => X"240F",
	003 => X"352B",
	004 => X"4533",
	005 => X"53D1",
	006 => X"60BB",
	007 => X"6BAD",
	008 => X"746D",
	009 => X"7ACF",
	010 => X"7EB1",
	011 => X"7FFF",
	012 => X"7EB1",
	013 => X"7ACF",
	014 => X"746D",
	015 => X"6BAD",
	016 => X"60BB",
	017 => X"53D1",
	018 => X"4533",
	019 => X"352B",
	020 => X"240F",
	021 => X"1237",
	022 => X"FFFD",
	023 => X"EDC6",
	024 => X"DBEE",
	025 => X"CAD2",
	026 => X"BACA",
	027 => X"AC2C",
	028 => X"9F42",
	029 => X"9450",
	030 => X"8B90",
	031 => X"852E",
	032 => X"814C",
	033 => X"7FFF",
	034 => X"814C",
	035 => X"852E",
	036 => X"8B90",
	037 => X"9450",
	038 => X"9F42",
	039 => X"AC2C",
	040 => X"BACA",
	041 => X"CAD2",
	042 => X"DBEE",
	043 => X"EDC6",
	044 => X"0000",
	045 => X"1237",
	046 => X"240F",
	047 => X"352B",
	048 => X"4533",
	049 => X"53D1",
	050 => X"60BB",
	051 => X"6BAD",
	052 => X"746D",
	053 => X"7ACF",
	054 => X"7EB1",
	055 => X"7FFF",
	056 => X"7EB1",
	057 => X"7ACF",
	058 => X"746D",
	059 => X"6BAD",
	060 => X"60BB",
	061 => X"53D1",
	062 => X"4533",
	063 => X"352B",
	064 => X"240F",
	065 => X"1237",
	066 => X"FFFD",
	067 => X"EDC6",
	068 => X"DBEE",
	069 => X"CAD2",
	070 => X"BACA",
	071 => X"AC2C",
	072 => X"9F42",
	073 => X"9450",
	074 => X"8B90",
	075 => X"852E",
	076 => X"814C",
	077 => X"7FFF",
	078 => X"814C",
	079 => X"852E",
	080 => X"8B90",
	081 => X"9450",
	082 => X"9F42",
	083 => X"AC2C",
	084 => X"BACA",
	085 => X"CAD2",
	086 => X"DBEE",
	087 => X"EDC6",
	088 => X"FFFD",
	089 => X"1237",
	090 => X"240F",
	091 => X"352B",
	092 => X"4533",
	093 => X"53D1",
	094 => X"60BB",
	095 => X"6BAD",
	096 => X"746D",
	097 => X"7ACF",
	098 => X"7EB1",
	099 => X"7FFF",
	100 => X"7EB1",
	101 => X"7ACF",
	102 => X"746D",
	103 => X"6BAD",
	104 => X"60BB",
	105 => X"53D1",
	106 => X"4533",
	107 => X"352B",
	108 => X"240F",
	109 => X"1237",
	110 => X"0000",
	111 => X"EDC6",
	112 => X"DBEE",
	113 => X"CAD2",
	114 => X"BACA",
	115 => X"AC2C",
	116 => X"9F42",
	117 => X"9450",
	118 => X"8B90",
	119 => X"852E",
	120 => X"814C",
	121 => X"7FFF",
	122 => X"814C",
	123 => X"852E",
	124 => X"8B90",
	125 => X"9450",
	126 => X"9F42",
	127 => X"AC2C",
	128 => X"BACA",
	129 => X"CAD2",
	130 => X"DBEE",
	131 => X"EDC6",
	132 => X"FFFD",
	133 => X"1237",
	134 => X"240F",
	135 => X"352B",
	136 => X"4533",
	137 => X"53D1",
	138 => X"60BB",
	139 => X"6BAD",
	140 => X"746D",
	141 => X"7ACF",
	142 => X"7EB1",
	143 => X"7FFF",
	144 => X"7EB1",
	145 => X"7ACF",
	146 => X"746D",
	147 => X"6BAD",
	148 => X"60BB",
	149 => X"53D1",
	150 => X"4533",
	151 => X"352B",
	152 => X"240F",
	153 => X"1237",
	154 => X"0000",
	155 => X"EDC6",
	156 => X"DBEE",
	157 => X"CAD2",
	158 => X"BACA",
	159 => X"AC2C",
	160 => X"9F42",
	161 => X"9450",
	162 => X"8B90",
	163 => X"852E",
	164 => X"814C",
	165 => X"7FFF",
	166 => X"814C",
	167 => X"852E",
	168 => X"8B90",
	169 => X"9450",
	170 => X"9F42",
	171 => X"AC2C",
	172 => X"BACA",
	173 => X"CAD2",
	174 => X"DBEE",
	175 => X"EDC6",
	176 => X"0000",
	177 => X"1237",
	178 => X"240F",
	179 => X"352B",
	180 => X"4533",
	181 => X"53D1",
	182 => X"60BB",
	183 => X"6BAD",
	184 => X"746D",
	185 => X"7ACF",
	186 => X"7EB1",
	187 => X"7FFF",
	188 => X"7EB1",
	189 => X"7ACF",
	190 => X"746D",
	191 => X"6BAD",
	192 => X"60BB",
	193 => X"53D1",
	194 => X"4533",
	195 => X"352B",
	196 => X"240F",
	197 => X"1237",
	198 => X"FFFD",
	199 => X"EDC6",
	200 => X"DBEE",
	201 => X"CAD2",
	202 => X"BACA",
	203 => X"AC2C",
	204 => X"9F42",
	205 => X"9450",
	206 => X"8B90",
	207 => X"852E",
	208 => X"814C",
	209 => X"7FFF",
	210 => X"814C",
	211 => X"852E",
	212 => X"8B90",
	213 => X"9450",
	214 => X"9F42",
	215 => X"AC2C",
	216 => X"BACA",
	217 => X"CAD2",
	218 => X"DBEE",
	219 => X"EDC6",
	220 => X"0000",
	221 => X"1237",
	222 => X"240F",
	223 => X"352B",
	224 => X"4533",
	225 => X"53D1",
	226 => X"60BB",
	227 => X"6BAD",
	228 => X"746D",
	229 => X"7ACF",
	230 => X"7EB1",
	231 => X"7FFF",
	232 => X"7EB1",
	233 => X"7ACF",
	234 => X"746D",
	235 => X"6BAD",
	236 => X"60BB",
	237 => X"53D1",
	238 => X"4533",
	239 => X"352B",
	240 => X"240F",
	241 => X"1237",
	242 => X"FFFD",
	243 => X"EDC6",
	244 => X"DBEE",
	245 => X"CAD2",
	246 => X"BACA",
	247 => X"AC2C",
	others => X"0000"
);

CONSTANT G5: hex := (
	000 => X"0000",
	001 => X"1313",
	002 => X"25BA",
	003 => X"3789",
	004 => X"481A",
	005 => X"570F",
	006 => X"6412",
	007 => X"6ED9",
	008 => X"7725",
	009 => X"7CC9",
	010 => X"7FA3",
	011 => X"7FA3",
	012 => X"7CC9",
	013 => X"7725",
	014 => X"6ED9",
	015 => X"6412",
	016 => X"570F",
	017 => X"481A",
	018 => X"3789",
	019 => X"25BA",
	020 => X"1313",
	021 => X"FFFD",
	022 => X"ECEA",
	023 => X"DA43",
	024 => X"C874",
	025 => X"B7E3",
	026 => X"A8EE",
	027 => X"9BEB",
	028 => X"9124",
	029 => X"88D8",
	030 => X"8334",
	031 => X"805A",
	032 => X"805A",
	033 => X"8334",
	034 => X"88D8",
	035 => X"9124",
	036 => X"9BEB",
	037 => X"A8EE",
	038 => X"B7E3",
	039 => X"C874",
	040 => X"DA43",
	041 => X"ECEA",
	042 => X"FFFD",
	043 => X"1313",
	044 => X"25BA",
	045 => X"3789",
	046 => X"481A",
	047 => X"570F",
	048 => X"6412",
	049 => X"6ED9",
	050 => X"7725",
	051 => X"7CC9",
	052 => X"7FA3",
	053 => X"7FA3",
	054 => X"7CC9",
	055 => X"7725",
	056 => X"6ED9",
	057 => X"6412",
	058 => X"570F",
	059 => X"481A",
	060 => X"3789",
	061 => X"25BA",
	062 => X"1313",
	063 => X"0000",
	064 => X"ECEA",
	065 => X"DA43",
	066 => X"C874",
	067 => X"B7E3",
	068 => X"A8EE",
	069 => X"9BEB",
	070 => X"9124",
	071 => X"88D8",
	072 => X"8334",
	073 => X"805A",
	074 => X"805A",
	075 => X"8334",
	076 => X"88D8",
	077 => X"9124",
	078 => X"9BEB",
	079 => X"A8EE",
	080 => X"B7E3",
	081 => X"C874",
	082 => X"DA43",
	083 => X"ECEA",
	084 => X"FFFD",
	085 => X"1313",
	086 => X"25BA",
	087 => X"3789",
	088 => X"481A",
	089 => X"570F",
	090 => X"6412",
	091 => X"6ED9",
	092 => X"7725",
	093 => X"7CC9",
	094 => X"7FA3",
	095 => X"7FA3",
	096 => X"7CC9",
	097 => X"7725",
	098 => X"6ED9",
	099 => X"6412",
	100 => X"570F",
	101 => X"481A",
	102 => X"3789",
	103 => X"25BA",
	104 => X"1313",
	105 => X"0000",
	106 => X"ECEA",
	107 => X"DA43",
	108 => X"C874",
	109 => X"B7E3",
	110 => X"A8EE",
	111 => X"9BEB",
	112 => X"9124",
	113 => X"88D8",
	114 => X"8334",
	115 => X"805A",
	116 => X"805A",
	117 => X"8334",
	118 => X"88D8",
	119 => X"9124",
	120 => X"9BEB",
	121 => X"A8EE",
	122 => X"B7E3",
	123 => X"C874",
	124 => X"DA43",
	125 => X"ECEA",
	126 => X"FFFD",
	127 => X"1313",
	128 => X"25BA",
	129 => X"3789",
	130 => X"481A",
	131 => X"570F",
	132 => X"6412",
	133 => X"6ED9",
	134 => X"7725",
	135 => X"7CC9",
	136 => X"7FA3",
	137 => X"7FA3",
	138 => X"7CC9",
	139 => X"7725",
	140 => X"6ED9",
	141 => X"6412",
	142 => X"570F",
	143 => X"481A",
	144 => X"3789",
	145 => X"25BA",
	146 => X"1313",
	147 => X"FFFD",
	148 => X"ECEA",
	149 => X"DA43",
	150 => X"C874",
	151 => X"B7E3",
	152 => X"A8EE",
	153 => X"9BEB",
	154 => X"9124",
	155 => X"88D8",
	156 => X"8334",
	157 => X"805A",
	158 => X"805A",
	159 => X"8334",
	160 => X"88D8",
	161 => X"9124",
	162 => X"9BEB",
	163 => X"A8EE",
	164 => X"B7E3",
	165 => X"C874",
	166 => X"DA43",
	167 => X"ECEA",
	168 => X"0000",
	169 => X"1313",
	170 => X"25BA",
	171 => X"3789",
	172 => X"481A",
	173 => X"570F",
	174 => X"6412",
	175 => X"6ED9",
	176 => X"7725",
	177 => X"7CC9",
	178 => X"7FA3",
	179 => X"7FA3",
	180 => X"7CC9",
	181 => X"7725",
	182 => X"6ED9",
	183 => X"6412",
	184 => X"570F",
	185 => X"481A",
	186 => X"3789",
	187 => X"25BA",
	188 => X"1313",
	189 => X"FFFD",
	190 => X"ECEA",
	191 => X"DA43",
	192 => X"C874",
	193 => X"B7E3",
	194 => X"A8EE",
	195 => X"9BEB",
	196 => X"9124",
	197 => X"88D8",
	198 => X"8334",
	199 => X"805A",
	200 => X"805A",
	201 => X"8334",
	202 => X"88D8",
	203 => X"9124",
	204 => X"9BEB",
	205 => X"A8EE",
	206 => X"B7E3",
	207 => X"C874",
	208 => X"DA43",
	209 => X"ECEA",
	210 => X"0000",
	211 => X"1313",
	212 => X"25BA",
	213 => X"3789",
	214 => X"481A",
	215 => X"570F",
	216 => X"6412",
	217 => X"6ED9",
	218 => X"7725",
	219 => X"7CC9",
	220 => X"7FA3",
	221 => X"7FA3",
	222 => X"7CC9",
	223 => X"7725",
	224 => X"6ED9",
	225 => X"6412",
	226 => X"570F",
	227 => X"481A",
	228 => X"3789",
	229 => X"25BA",
	230 => X"1313",
	231 => X"FFFD",
	232 => X"ECEA",
	233 => X"DA43",
	234 => X"C874",
	235 => X"B7E3",
	236 => X"A8EE",
	237 => X"9BEB",
	238 => X"9124",
	239 => X"88D8",
	240 => X"8334",
	241 => X"805A",
	242 => X"805A",
	243 => X"8334",
	244 => X"88D8",
	245 => X"9124",
	246 => X"9BEB",
	247 => X"A8EE",
	others => X"0000"
);

CONSTANT GS5: hex := (
	000 => X"0000",
	001 => X"1488",
	002 => X"2888",
	003 => X"3B7B",
	004 => X"4CE4",
	005 => X"5C4F",
	006 => X"6956",
	007 => X"73A3",
	008 => X"7AF1",
	009 => X"7F10",
	010 => X"7FE4",
	011 => X"7D68",
	012 => X"77AD",
	013 => X"6ED9",
	014 => X"6325",
	015 => X"54E0",
	016 => X"4468",
	017 => X"322B",
	018 => X"1EA1",
	019 => X"0A4C",
	020 => X"F5B1",
	021 => X"E15C",
	022 => X"CDD2",
	023 => X"BB95",
	024 => X"AB1D",
	025 => X"9CD8",
	026 => X"9124",
	027 => X"8850",
	028 => X"8295",
	029 => X"8019",
	030 => X"80ED",
	031 => X"850C",
	032 => X"8C5A",
	033 => X"96A7",
	034 => X"A3AE",
	035 => X"B319",
	036 => X"C482",
	037 => X"D775",
	038 => X"EB75",
	039 => X"FFFD",
	040 => X"1488",
	041 => X"2888",
	042 => X"3B7B",
	043 => X"4CE4",
	044 => X"5C4F",
	045 => X"6956",
	046 => X"73A3",
	047 => X"7AF1",
	048 => X"7F10",
	049 => X"7FE4",
	050 => X"7D68",
	051 => X"77AD",
	052 => X"6ED9",
	053 => X"6325",
	054 => X"54E0",
	055 => X"4468",
	056 => X"322B",
	057 => X"1EA1",
	058 => X"0A4C",
	059 => X"F5B1",
	060 => X"E15C",
	061 => X"CDD2",
	062 => X"BB95",
	063 => X"AB1D",
	064 => X"9CD8",
	065 => X"9124",
	066 => X"8850",
	067 => X"8295",
	068 => X"8019",
	069 => X"80ED",
	070 => X"850C",
	071 => X"8C5A",
	072 => X"96A7",
	073 => X"A3AE",
	074 => X"B319",
	075 => X"C482",
	076 => X"D775",
	077 => X"EB75",
	078 => X"0000",
	079 => X"1488",
	080 => X"2888",
	081 => X"3B7B",
	082 => X"4CE4",
	083 => X"5C4F",
	084 => X"6956",
	085 => X"73A3",
	086 => X"7AF1",
	087 => X"7F10",
	088 => X"7FE4",
	089 => X"7D68",
	090 => X"77AD",
	091 => X"6ED9",
	092 => X"6325",
	093 => X"54E0",
	094 => X"4468",
	095 => X"322B",
	096 => X"1EA1",
	097 => X"0A4C",
	098 => X"F5B1",
	099 => X"E15C",
	100 => X"CDD2",
	101 => X"BB95",
	102 => X"AB1D",
	103 => X"9CD8",
	104 => X"9124",
	105 => X"8850",
	106 => X"8295",
	107 => X"8019",
	108 => X"80ED",
	109 => X"850C",
	110 => X"8C5A",
	111 => X"96A7",
	112 => X"A3AE",
	113 => X"B319",
	114 => X"C482",
	115 => X"D775",
	116 => X"EB75",
	117 => X"0000",
	118 => X"1488",
	119 => X"2888",
	120 => X"3B7B",
	121 => X"4CE4",
	122 => X"5C4F",
	123 => X"6956",
	124 => X"73A3",
	125 => X"7AF1",
	126 => X"7F10",
	127 => X"7FE4",
	128 => X"7D68",
	129 => X"77AD",
	130 => X"6ED9",
	131 => X"6325",
	132 => X"54E0",
	133 => X"4468",
	134 => X"322B",
	135 => X"1EA1",
	136 => X"0A4C",
	137 => X"F5B1",
	138 => X"E15C",
	139 => X"CDD2",
	140 => X"BB95",
	141 => X"AB1D",
	142 => X"9CD8",
	143 => X"9124",
	144 => X"8850",
	145 => X"8295",
	146 => X"8019",
	147 => X"80ED",
	148 => X"850C",
	149 => X"8C5A",
	150 => X"96A7",
	151 => X"A3AE",
	152 => X"B319",
	153 => X"C482",
	154 => X"D775",
	155 => X"EB75",
	156 => X"0000",
	157 => X"1488",
	158 => X"2888",
	159 => X"3B7B",
	160 => X"4CE4",
	161 => X"5C4F",
	162 => X"6956",
	163 => X"73A3",
	164 => X"7AF1",
	165 => X"7F10",
	166 => X"7FE4",
	167 => X"7D68",
	168 => X"77AD",
	169 => X"6ED9",
	170 => X"6325",
	171 => X"54E0",
	172 => X"4468",
	173 => X"322B",
	174 => X"1EA1",
	175 => X"0A4C",
	176 => X"F5B1",
	177 => X"E15C",
	178 => X"CDD2",
	179 => X"BB95",
	180 => X"AB1D",
	181 => X"9CD8",
	182 => X"9124",
	183 => X"8850",
	184 => X"8295",
	185 => X"8019",
	186 => X"80ED",
	187 => X"850C",
	188 => X"8C5A",
	189 => X"96A7",
	190 => X"A3AE",
	191 => X"B319",
	192 => X"C482",
	193 => X"D775",
	194 => X"EB75",
	195 => X"0000",
	196 => X"1488",
	197 => X"2888",
	198 => X"3B7B",
	199 => X"4CE4",
	200 => X"5C4F",
	201 => X"6956",
	202 => X"73A3",
	203 => X"7AF1",
	204 => X"7F10",
	205 => X"7FE4",
	206 => X"7D68",
	207 => X"77AD",
	208 => X"6ED9",
	209 => X"6325",
	210 => X"54E0",
	211 => X"4468",
	212 => X"322B",
	213 => X"1EA1",
	214 => X"0A4C",
	215 => X"F5B1",
	216 => X"E15C",
	217 => X"CDD2",
	218 => X"BB95",
	219 => X"AB1D",
	220 => X"9CD8",
	221 => X"9124",
	222 => X"8850",
	223 => X"8295",
	224 => X"8019",
	225 => X"80ED",
	226 => X"850C",
	227 => X"8C5A",
	228 => X"96A7",
	229 => X"A3AE",
	230 => X"B319",
	231 => X"C482",
	232 => X"D775",
	233 => X"EB75",
	234 => X"0000",
	235 => X"1488",
	236 => X"2888",
	237 => X"3B7B",
	238 => X"4CE4",
	239 => X"5C4F",
	240 => X"6956",
	241 => X"73A3",
	242 => X"7AF1",
	243 => X"7F10",
	244 => X"7FE4",
	245 => X"7D68",
	246 => X"77AD",
	247 => X"6ED9",
	others => X"0000"
);

CONSTANT A5: hex := (
	000 => X"0000",
	001 => X"15A1",
	002 => X"2AA3",
	003 => X"3E6C",
	004 => X"5068",
	005 => X"6015",
	006 => X"6CFE",
	007 => X"76C4",
	008 => X"7D1F",
	009 => X"7FE1",
	010 => X"7EF5",
	011 => X"7A62",
	012 => X"724A",
	013 => X"66E8",
	014 => X"5890",
	015 => X"47AC",
	016 => X"34B8",
	017 => X"2040",
	018 => X"0ADA",
	019 => X"F523",
	020 => X"DFBD",
	021 => X"CB45",
	022 => X"B851",
	023 => X"A76D",
	024 => X"9915",
	025 => X"8DB3",
	026 => X"859B",
	027 => X"8108",
	028 => X"801C",
	029 => X"82DE",
	030 => X"8939",
	031 => X"92FF",
	032 => X"9FE8",
	033 => X"AF95",
	034 => X"C191",
	035 => X"D55A",
	036 => X"EA5C",
	037 => X"0000",
	038 => X"15A1",
	039 => X"2AA3",
	040 => X"3E6C",
	041 => X"5068",
	042 => X"6015",
	043 => X"6CFE",
	044 => X"76C4",
	045 => X"7D1F",
	046 => X"7FE1",
	047 => X"7EF5",
	048 => X"7A62",
	049 => X"724A",
	050 => X"66E8",
	051 => X"5890",
	052 => X"47AC",
	053 => X"34B8",
	054 => X"2040",
	055 => X"0ADA",
	056 => X"F523",
	057 => X"DFBD",
	058 => X"CB45",
	059 => X"B851",
	060 => X"A76D",
	061 => X"9915",
	062 => X"8DB3",
	063 => X"859B",
	064 => X"8108",
	065 => X"801C",
	066 => X"82DE",
	067 => X"8939",
	068 => X"92FF",
	069 => X"9FE8",
	070 => X"AF95",
	071 => X"C191",
	072 => X"D55A",
	073 => X"EA5C",
	074 => X"FFFD",
	075 => X"15A1",
	076 => X"2AA3",
	077 => X"3E6C",
	078 => X"5068",
	079 => X"6015",
	080 => X"6CFE",
	081 => X"76C4",
	082 => X"7D1F",
	083 => X"7FE1",
	084 => X"7EF5",
	085 => X"7A62",
	086 => X"724A",
	087 => X"66E8",
	088 => X"5890",
	089 => X"47AC",
	090 => X"34B8",
	091 => X"2040",
	092 => X"0ADA",
	093 => X"F523",
	094 => X"DFBD",
	095 => X"CB45",
	096 => X"B851",
	097 => X"A76D",
	098 => X"9915",
	099 => X"8DB3",
	100 => X"859B",
	101 => X"8108",
	102 => X"801C",
	103 => X"82DE",
	104 => X"8939",
	105 => X"92FF",
	106 => X"9FE8",
	107 => X"AF95",
	108 => X"C191",
	109 => X"D55A",
	110 => X"EA5C",
	111 => X"FFFD",
	112 => X"15A1",
	113 => X"2AA3",
	114 => X"3E6C",
	115 => X"5068",
	116 => X"6015",
	117 => X"6CFE",
	118 => X"76C4",
	119 => X"7D1F",
	120 => X"7FE1",
	121 => X"7EF5",
	122 => X"7A62",
	123 => X"724A",
	124 => X"66E8",
	125 => X"5890",
	126 => X"47AC",
	127 => X"34B8",
	128 => X"2040",
	129 => X"0ADA",
	130 => X"F523",
	131 => X"DFBD",
	132 => X"CB45",
	133 => X"B851",
	134 => X"A76D",
	135 => X"9915",
	136 => X"8DB3",
	137 => X"859B",
	138 => X"8108",
	139 => X"801C",
	140 => X"82DE",
	141 => X"8939",
	142 => X"92FF",
	143 => X"9FE8",
	144 => X"AF95",
	145 => X"C191",
	146 => X"D55A",
	147 => X"EA5C",
	148 => X"0000",
	149 => X"15A1",
	150 => X"2AA3",
	151 => X"3E6C",
	152 => X"5068",
	153 => X"6015",
	154 => X"6CFE",
	155 => X"76C4",
	156 => X"7D1F",
	157 => X"7FE1",
	158 => X"7EF5",
	159 => X"7A62",
	160 => X"724A",
	161 => X"66E8",
	162 => X"5890",
	163 => X"47AC",
	164 => X"34B8",
	165 => X"2040",
	166 => X"0ADA",
	167 => X"F523",
	168 => X"DFBD",
	169 => X"CB45",
	170 => X"B851",
	171 => X"A76D",
	172 => X"9915",
	173 => X"8DB3",
	174 => X"859B",
	175 => X"8108",
	176 => X"801C",
	177 => X"82DE",
	178 => X"8939",
	179 => X"92FF",
	180 => X"9FE8",
	181 => X"AF95",
	182 => X"C191",
	183 => X"D55A",
	184 => X"EA5C",
	185 => X"0000",
	186 => X"15A1",
	187 => X"2AA3",
	188 => X"3E6C",
	189 => X"5068",
	190 => X"6015",
	191 => X"6CFE",
	192 => X"76C4",
	193 => X"7D1F",
	194 => X"7FE1",
	195 => X"7EF5",
	196 => X"7A62",
	197 => X"724A",
	198 => X"66E8",
	199 => X"5890",
	200 => X"47AC",
	201 => X"34B8",
	202 => X"2040",
	203 => X"0ADA",
	204 => X"F523",
	205 => X"DFBD",
	206 => X"CB45",
	207 => X"B851",
	208 => X"A76D",
	209 => X"9915",
	210 => X"8DB3",
	211 => X"859B",
	212 => X"8108",
	213 => X"801C",
	214 => X"82DE",
	215 => X"8939",
	216 => X"92FF",
	217 => X"9FE8",
	218 => X"AF95",
	219 => X"C191",
	220 => X"D55A",
	221 => X"EA5C",
	222 => X"0000",
	223 => X"15A1",
	224 => X"2AA3",
	225 => X"3E6C",
	226 => X"5068",
	227 => X"6015",
	228 => X"6CFE",
	229 => X"76C4",
	230 => X"7D1F",
	231 => X"7FE1",
	232 => X"7EF5",
	233 => X"7A62",
	234 => X"724A",
	235 => X"66E8",
	236 => X"5890",
	237 => X"47AC",
	238 => X"34B8",
	239 => X"2040",
	240 => X"0ADA",
	241 => X"F523",
	242 => X"DFBD",
	243 => X"CB45",
	244 => X"B851",
	245 => X"A76D",
	246 => X"9915",
	247 => X"8DB3",
	others => X"0000"
);

CONSTANT AS5: hex := (
	000 => X"0000",
	001 => X"16DA",
	002 => X"2CF9",
	003 => X"41A6",
	004 => X"5436",
	005 => X"6412",
	006 => X"70B6",
	007 => X"79BB",
	008 => X"7ED6",
	009 => X"7FDE",
	010 => X"7CC9",
	011 => X"75B2",
	012 => X"6AD2",
	013 => X"5C83",
	014 => X"4B3B",
	015 => X"3789",
	016 => X"220D",
	017 => X"0B79",
	018 => X"F484",
	019 => X"DDF0",
	020 => X"C874",
	021 => X"B4C2",
	022 => X"A37A",
	023 => X"952B",
	024 => X"8A4B",
	025 => X"8334",
	026 => X"801F",
	027 => X"8127",
	028 => X"8642",
	029 => X"8F47",
	030 => X"9BEB",
	031 => X"ABC7",
	032 => X"BE57",
	033 => X"D304",
	034 => X"E923",
	035 => X"FFFD",
	036 => X"16DA",
	037 => X"2CF9",
	038 => X"41A6",
	039 => X"5436",
	040 => X"6412",
	041 => X"70B6",
	042 => X"79BB",
	043 => X"7ED6",
	044 => X"7FDE",
	045 => X"7CC9",
	046 => X"75B2",
	047 => X"6AD2",
	048 => X"5C83",
	049 => X"4B3B",
	050 => X"3789",
	051 => X"220D",
	052 => X"0B79",
	053 => X"F484",
	054 => X"DDF0",
	055 => X"C874",
	056 => X"B4C2",
	057 => X"A37A",
	058 => X"952B",
	059 => X"8A4B",
	060 => X"8334",
	061 => X"801F",
	062 => X"8127",
	063 => X"8642",
	064 => X"8F47",
	065 => X"9BEB",
	066 => X"ABC7",
	067 => X"BE57",
	068 => X"D304",
	069 => X"E923",
	070 => X"0000",
	071 => X"16DA",
	072 => X"2CF9",
	073 => X"41A6",
	074 => X"5436",
	075 => X"6412",
	076 => X"70B6",
	077 => X"79BB",
	078 => X"7ED6",
	079 => X"7FDE",
	080 => X"7CC9",
	081 => X"75B2",
	082 => X"6AD2",
	083 => X"5C83",
	084 => X"4B3B",
	085 => X"3789",
	086 => X"220D",
	087 => X"0B79",
	088 => X"F484",
	089 => X"DDF0",
	090 => X"C874",
	091 => X"B4C2",
	092 => X"A37A",
	093 => X"952B",
	094 => X"8A4B",
	095 => X"8334",
	096 => X"801F",
	097 => X"8127",
	098 => X"8642",
	099 => X"8F47",
	100 => X"9BEB",
	101 => X"ABC7",
	102 => X"BE57",
	103 => X"D304",
	104 => X"E923",
	105 => X"0000",
	106 => X"16DA",
	107 => X"2CF9",
	108 => X"41A6",
	109 => X"5436",
	110 => X"6412",
	111 => X"70B6",
	112 => X"79BB",
	113 => X"7ED6",
	114 => X"7FDE",
	115 => X"7CC9",
	116 => X"75B2",
	117 => X"6AD2",
	118 => X"5C83",
	119 => X"4B3B",
	120 => X"3789",
	121 => X"220D",
	122 => X"0B79",
	123 => X"F484",
	124 => X"DDF0",
	125 => X"C874",
	126 => X"B4C2",
	127 => X"A37A",
	128 => X"952B",
	129 => X"8A4B",
	130 => X"8334",
	131 => X"801F",
	132 => X"8127",
	133 => X"8642",
	134 => X"8F47",
	135 => X"9BEB",
	136 => X"ABC7",
	137 => X"BE57",
	138 => X"D304",
	139 => X"E923",
	140 => X"FFFD",
	141 => X"16DA",
	142 => X"2CF9",
	143 => X"41A6",
	144 => X"5436",
	145 => X"6412",
	146 => X"70B6",
	147 => X"79BB",
	148 => X"7ED6",
	149 => X"7FDE",
	150 => X"7CC9",
	151 => X"75B2",
	152 => X"6AD2",
	153 => X"5C83",
	154 => X"4B3B",
	155 => X"3789",
	156 => X"220D",
	157 => X"0B79",
	158 => X"F484",
	159 => X"DDF0",
	160 => X"C874",
	161 => X"B4C2",
	162 => X"A37A",
	163 => X"952B",
	164 => X"8A4B",
	165 => X"8334",
	166 => X"801F",
	167 => X"8127",
	168 => X"8642",
	169 => X"8F47",
	170 => X"9BEB",
	171 => X"ABC7",
	172 => X"BE57",
	173 => X"D304",
	174 => X"E923",
	175 => X"FFFD",
	176 => X"16DA",
	177 => X"2CF9",
	178 => X"41A6",
	179 => X"5436",
	180 => X"6412",
	181 => X"70B6",
	182 => X"79BB",
	183 => X"7ED6",
	184 => X"7FDE",
	185 => X"7CC9",
	186 => X"75B2",
	187 => X"6AD2",
	188 => X"5C83",
	189 => X"4B3B",
	190 => X"3789",
	191 => X"220D",
	192 => X"0B79",
	193 => X"F484",
	194 => X"DDF0",
	195 => X"C874",
	196 => X"B4C2",
	197 => X"A37A",
	198 => X"952B",
	199 => X"8A4B",
	200 => X"8334",
	201 => X"801F",
	202 => X"8127",
	203 => X"8642",
	204 => X"8F47",
	205 => X"9BEB",
	206 => X"ABC7",
	207 => X"BE57",
	208 => X"D304",
	209 => X"E923",
	210 => X"FFFD",
	211 => X"16DA",
	212 => X"2CF9",
	213 => X"41A6",
	214 => X"5436",
	215 => X"6412",
	216 => X"70B6",
	217 => X"79BB",
	218 => X"7ED6",
	219 => X"7FDE",
	220 => X"7CC9",
	221 => X"75B2",
	222 => X"6AD2",
	223 => X"5C83",
	224 => X"4B3B",
	225 => X"3789",
	226 => X"220D",
	227 => X"0B79",
	228 => X"F484",
	229 => X"DDF0",
	230 => X"C874",
	231 => X"B4C2",
	232 => X"A37A",
	233 => X"952B",
	234 => X"8A4B",
	235 => X"8334",
	236 => X"801F",
	237 => X"8127",
	238 => X"8642",
	239 => X"8F47",
	240 => X"9BEB",
	241 => X"ABC7",
	242 => X"BE57",
	243 => X"D304",
	244 => X"E923",
	245 => X"FFFD",
	246 => X"16DA",
	247 => X"2CF9",
	others => X"0000"
);

CONSTANT B5: hex := (
	000 => X"0000",
	001 => X"1839",
	002 => X"2F92",
	003 => X"4533",
	004 => X"5853",
	005 => X"6843",
	006 => X"746D",
	007 => X"7C63",
	008 => X"7FD9",
	009 => X"7EB1",
	010 => X"78F4",
	011 => X"6ED9",
	012 => X"60BB",
	013 => X"4F1F",
	014 => X"3AA6",
	015 => X"240F",
	016 => X"0C2A",
	017 => X"F3D3",
	018 => X"DBEE",
	019 => X"C557",
	020 => X"B0DE",
	021 => X"9F42",
	022 => X"9124",
	023 => X"8709",
	024 => X"814C",
	025 => X"8024",
	026 => X"839A",
	027 => X"8B90",
	028 => X"97BA",
	029 => X"A7AA",
	030 => X"BACA",
	031 => X"D06B",
	032 => X"E7C4",
	033 => X"0000",
	034 => X"1839",
	035 => X"2F92",
	036 => X"4533",
	037 => X"5853",
	038 => X"6843",
	039 => X"746D",
	040 => X"7C63",
	041 => X"7FD9",
	042 => X"7EB1",
	043 => X"78F4",
	044 => X"6ED9",
	045 => X"60BB",
	046 => X"4F1F",
	047 => X"3AA6",
	048 => X"240F",
	049 => X"0C2A",
	050 => X"F3D3",
	051 => X"DBEE",
	052 => X"C557",
	053 => X"B0DE",
	054 => X"9F42",
	055 => X"9124",
	056 => X"8709",
	057 => X"814C",
	058 => X"8024",
	059 => X"839A",
	060 => X"8B90",
	061 => X"97BA",
	062 => X"A7AA",
	063 => X"BACA",
	064 => X"D06B",
	065 => X"E7C4",
	066 => X"FFFD",
	067 => X"1839",
	068 => X"2F92",
	069 => X"4533",
	070 => X"5853",
	071 => X"6843",
	072 => X"746D",
	073 => X"7C63",
	074 => X"7FD9",
	075 => X"7EB1",
	076 => X"78F4",
	077 => X"6ED9",
	078 => X"60BB",
	079 => X"4F1F",
	080 => X"3AA6",
	081 => X"240F",
	082 => X"0C2A",
	083 => X"F3D3",
	084 => X"DBEE",
	085 => X"C557",
	086 => X"B0DE",
	087 => X"9F42",
	088 => X"9124",
	089 => X"8709",
	090 => X"814C",
	091 => X"8024",
	092 => X"839A",
	093 => X"8B90",
	094 => X"97BA",
	095 => X"A7AA",
	096 => X"BACA",
	097 => X"D06B",
	098 => X"E7C4",
	099 => X"FFFD",
	100 => X"1839",
	101 => X"2F92",
	102 => X"4533",
	103 => X"5853",
	104 => X"6843",
	105 => X"746D",
	106 => X"7C63",
	107 => X"7FD9",
	108 => X"7EB1",
	109 => X"78F4",
	110 => X"6ED9",
	111 => X"60BB",
	112 => X"4F1F",
	113 => X"3AA6",
	114 => X"240F",
	115 => X"0C2A",
	116 => X"F3D3",
	117 => X"DBEE",
	118 => X"C557",
	119 => X"B0DE",
	120 => X"9F42",
	121 => X"9124",
	122 => X"8709",
	123 => X"814C",
	124 => X"8024",
	125 => X"839A",
	126 => X"8B90",
	127 => X"97BA",
	128 => X"A7AA",
	129 => X"BACA",
	130 => X"D06B",
	131 => X"E7C4",
	132 => X"0000",
	133 => X"1839",
	134 => X"2F92",
	135 => X"4533",
	136 => X"5853",
	137 => X"6843",
	138 => X"746D",
	139 => X"7C63",
	140 => X"7FD9",
	141 => X"7EB1",
	142 => X"78F4",
	143 => X"6ED9",
	144 => X"60BB",
	145 => X"4F1F",
	146 => X"3AA6",
	147 => X"240F",
	148 => X"0C2A",
	149 => X"F3D3",
	150 => X"DBEE",
	151 => X"C557",
	152 => X"B0DE",
	153 => X"9F42",
	154 => X"9124",
	155 => X"8709",
	156 => X"814C",
	157 => X"8024",
	158 => X"839A",
	159 => X"8B90",
	160 => X"97BA",
	161 => X"A7AA",
	162 => X"BACA",
	163 => X"D06B",
	164 => X"E7C4",
	165 => X"0000",
	166 => X"1839",
	167 => X"2F92",
	168 => X"4533",
	169 => X"5853",
	170 => X"6843",
	171 => X"746D",
	172 => X"7C63",
	173 => X"7FD9",
	174 => X"7EB1",
	175 => X"78F4",
	176 => X"6ED9",
	177 => X"60BB",
	178 => X"4F1F",
	179 => X"3AA6",
	180 => X"240F",
	181 => X"0C2A",
	182 => X"F3D3",
	183 => X"DBEE",
	184 => X"C557",
	185 => X"B0DE",
	186 => X"9F42",
	187 => X"9124",
	188 => X"8709",
	189 => X"814C",
	190 => X"8024",
	191 => X"839A",
	192 => X"8B90",
	193 => X"97BA",
	194 => X"A7AA",
	195 => X"BACA",
	196 => X"D06B",
	197 => X"E7C4",
	198 => X"0000",
	199 => X"1839",
	200 => X"2F92",
	201 => X"4533",
	202 => X"5853",
	203 => X"6843",
	204 => X"746D",
	205 => X"7C63",
	206 => X"7FD9",
	207 => X"7EB1",
	208 => X"78F4",
	209 => X"6ED9",
	210 => X"60BB",
	211 => X"4F1F",
	212 => X"3AA6",
	213 => X"240F",
	214 => X"0C2A",
	215 => X"F3D3",
	216 => X"DBEE",
	217 => X"C557",
	218 => X"B0DE",
	219 => X"9F42",
	220 => X"9124",
	221 => X"8709",
	222 => X"814C",
	223 => X"8024",
	224 => X"839A",
	225 => X"8B90",
	226 => X"97BA",
	227 => X"A7AA",
	228 => X"BACA",
	229 => X"D06B",
	230 => X"E7C4",
	231 => X"0000",
	232 => X"1839",
	233 => X"2F92",
	234 => X"4533",
	235 => X"5853",
	236 => X"6843",
	237 => X"746D",
	238 => X"7C63",
	239 => X"7FD9",
	240 => X"7EB1",
	241 => X"78F4",
	242 => X"6ED9",
	243 => X"60BB",
	244 => X"4F1F",
	245 => X"3AA6",
	246 => X"240F",
	247 => X"0C2A",
	others => X"0000"
);

CONSTANT C6: hex := (
	000 => X"0000",
	001 => X"19C3",
	002 => X"3279",
	003 => X"491E",
	004 => X"5CC5",
	005 => X"6C9F",
	006 => X"7807",
	007 => X"7E85",
	008 => X"7FD4",
	009 => X"7BE8",
	010 => X"72EA",
	011 => X"6537",
	012 => X"535F",
	013 => X"3E1D",
	014 => X"2651",
	015 => X"0CF2",
	016 => X"F30B",
	017 => X"D9AC",
	018 => X"C1E0",
	019 => X"AC9E",
	020 => X"9AC6",
	021 => X"8D13",
	022 => X"8415",
	023 => X"8029",
	024 => X"8178",
	025 => X"87F6",
	026 => X"935E",
	027 => X"A338",
	028 => X"B6DF",
	029 => X"CD84",
	030 => X"E63A",
	031 => X"0000",
	032 => X"19C3",
	033 => X"3279",
	034 => X"491E",
	035 => X"5CC5",
	036 => X"6C9F",
	037 => X"7807",
	038 => X"7E85",
	039 => X"7FD4",
	040 => X"7BE8",
	041 => X"72EA",
	042 => X"6537",
	043 => X"535F",
	044 => X"3E1D",
	045 => X"2651",
	046 => X"0CF2",
	047 => X"F30B",
	048 => X"D9AC",
	049 => X"C1E0",
	050 => X"AC9E",
	051 => X"9AC6",
	052 => X"8D13",
	053 => X"8415",
	054 => X"8029",
	055 => X"8178",
	056 => X"87F6",
	057 => X"935E",
	058 => X"A338",
	059 => X"B6DF",
	060 => X"CD84",
	061 => X"E63A",
	062 => X"0000",
	063 => X"19C3",
	064 => X"3279",
	065 => X"491E",
	066 => X"5CC5",
	067 => X"6C9F",
	068 => X"7807",
	069 => X"7E85",
	070 => X"7FD4",
	071 => X"7BE8",
	072 => X"72EA",
	073 => X"6537",
	074 => X"535F",
	075 => X"3E1D",
	076 => X"2651",
	077 => X"0CF2",
	078 => X"F30B",
	079 => X"D9AC",
	080 => X"C1E0",
	081 => X"AC9E",
	082 => X"9AC6",
	083 => X"8D13",
	084 => X"8415",
	085 => X"8029",
	086 => X"8178",
	087 => X"87F6",
	088 => X"935E",
	089 => X"A338",
	090 => X"B6DF",
	091 => X"CD84",
	092 => X"E63A",
	093 => X"0000",
	094 => X"19C3",
	095 => X"3279",
	096 => X"491E",
	097 => X"5CC5",
	098 => X"6C9F",
	099 => X"7807",
	100 => X"7E85",
	101 => X"7FD4",
	102 => X"7BE8",
	103 => X"72EA",
	104 => X"6537",
	105 => X"535F",
	106 => X"3E1D",
	107 => X"2651",
	108 => X"0CF2",
	109 => X"F30B",
	110 => X"D9AC",
	111 => X"C1E0",
	112 => X"AC9E",
	113 => X"9AC6",
	114 => X"8D13",
	115 => X"8415",
	116 => X"8029",
	117 => X"8178",
	118 => X"87F6",
	119 => X"935E",
	120 => X"A338",
	121 => X"B6DF",
	122 => X"CD84",
	123 => X"E63A",
	124 => X"FFFD",
	125 => X"19C3",
	126 => X"3279",
	127 => X"491E",
	128 => X"5CC5",
	129 => X"6C9F",
	130 => X"7807",
	131 => X"7E85",
	132 => X"7FD4",
	133 => X"7BE8",
	134 => X"72EA",
	135 => X"6537",
	136 => X"535F",
	137 => X"3E1D",
	138 => X"2651",
	139 => X"0CF2",
	140 => X"F30B",
	141 => X"D9AC",
	142 => X"C1E0",
	143 => X"AC9E",
	144 => X"9AC6",
	145 => X"8D13",
	146 => X"8415",
	147 => X"8029",
	148 => X"8178",
	149 => X"87F6",
	150 => X"935E",
	151 => X"A338",
	152 => X"B6DF",
	153 => X"CD84",
	154 => X"E63A",
	155 => X"FFFD",
	156 => X"19C3",
	157 => X"3279",
	158 => X"491E",
	159 => X"5CC5",
	160 => X"6C9F",
	161 => X"7807",
	162 => X"7E85",
	163 => X"7FD4",
	164 => X"7BE8",
	165 => X"72EA",
	166 => X"6537",
	167 => X"535F",
	168 => X"3E1D",
	169 => X"2651",
	170 => X"0CF2",
	171 => X"F30B",
	172 => X"D9AC",
	173 => X"C1E0",
	174 => X"AC9E",
	175 => X"9AC6",
	176 => X"8D13",
	177 => X"8415",
	178 => X"8029",
	179 => X"8178",
	180 => X"87F6",
	181 => X"935E",
	182 => X"A338",
	183 => X"B6DF",
	184 => X"CD84",
	185 => X"E63A",
	186 => X"FFFD",
	187 => X"19C3",
	188 => X"3279",
	189 => X"491E",
	190 => X"5CC5",
	191 => X"6C9F",
	192 => X"7807",
	193 => X"7E85",
	194 => X"7FD4",
	195 => X"7BE8",
	196 => X"72EA",
	197 => X"6537",
	198 => X"535F",
	199 => X"3E1D",
	200 => X"2651",
	201 => X"0CF2",
	202 => X"F30B",
	203 => X"D9AC",
	204 => X"C1E0",
	205 => X"AC9E",
	206 => X"9AC6",
	207 => X"8D13",
	208 => X"8415",
	209 => X"8029",
	210 => X"8178",
	211 => X"87F6",
	212 => X"935E",
	213 => X"A338",
	214 => X"B6DF",
	215 => X"CD84",
	216 => X"E63A",
	217 => X"FFFD",
	218 => X"19C3",
	219 => X"3279",
	220 => X"491E",
	221 => X"5CC5",
	222 => X"6C9F",
	223 => X"7807",
	224 => X"7E85",
	225 => X"7FD4",
	226 => X"7BE8",
	227 => X"72EA",
	228 => X"6537",
	229 => X"535F",
	230 => X"3E1D",
	231 => X"2651",
	232 => X"0CF2",
	233 => X"F30B",
	234 => X"D9AC",
	235 => X"C1E0",
	236 => X"AC9E",
	237 => X"9AC6",
	238 => X"8D13",
	239 => X"8415",
	240 => X"8029",
	241 => X"8178",
	242 => X"87F6",
	243 => X"935E",
	244 => X"A338",
	245 => X"B6DF",
	246 => X"CD84",
	247 => X"E63A",
	others => X"0000"
);

CONSTANT CS6: hex := (
	000 => X"0000",
	001 => X"1B83",
	002 => X"35BE",
	003 => X"4D75",
	004 => X"618D",
	005 => X"7116",
	006 => X"7B54",
	007 => X"7FCE",
	008 => X"7E4F",
	009 => X"76E7",
	010 => X"69F0",
	011 => X"5805",
	012 => X"41FD",
	013 => X"28DE",
	014 => X"0DD6",
	015 => X"F227",
	016 => X"D71F",
	017 => X"BE00",
	018 => X"A7F8",
	019 => X"960D",
	020 => X"8916",
	021 => X"81AE",
	022 => X"802F",
	023 => X"84A9",
	024 => X"8EE7",
	025 => X"9E70",
	026 => X"B288",
	027 => X"CA3F",
	028 => X"E47A",
	029 => X"FFFD",
	030 => X"1B83",
	031 => X"35BE",
	032 => X"4D75",
	033 => X"618D",
	034 => X"7116",
	035 => X"7B54",
	036 => X"7FCE",
	037 => X"7E4F",
	038 => X"76E7",
	039 => X"69F0",
	040 => X"5805",
	041 => X"41FD",
	042 => X"28DE",
	043 => X"0DD6",
	044 => X"F227",
	045 => X"D71F",
	046 => X"BE00",
	047 => X"A7F8",
	048 => X"960D",
	049 => X"8916",
	050 => X"81AE",
	051 => X"802F",
	052 => X"84A9",
	053 => X"8EE7",
	054 => X"9E70",
	055 => X"B288",
	056 => X"CA3F",
	057 => X"E47A",
	058 => X"FFFD",
	059 => X"1B83",
	060 => X"35BE",
	061 => X"4D75",
	062 => X"618D",
	063 => X"7116",
	064 => X"7B54",
	065 => X"7FCE",
	066 => X"7E4F",
	067 => X"76E7",
	068 => X"69F0",
	069 => X"5805",
	070 => X"41FD",
	071 => X"28DE",
	072 => X"0DD6",
	073 => X"F227",
	074 => X"D71F",
	075 => X"BE00",
	076 => X"A7F8",
	077 => X"960D",
	078 => X"8916",
	079 => X"81AE",
	080 => X"802F",
	081 => X"84A9",
	082 => X"8EE7",
	083 => X"9E70",
	084 => X"B288",
	085 => X"CA3F",
	086 => X"E47A",
	087 => X"FFFD",
	088 => X"1B83",
	089 => X"35BE",
	090 => X"4D75",
	091 => X"618D",
	092 => X"7116",
	093 => X"7B54",
	094 => X"7FCE",
	095 => X"7E4F",
	096 => X"76E7",
	097 => X"69F0",
	098 => X"5805",
	099 => X"41FD",
	100 => X"28DE",
	101 => X"0DD6",
	102 => X"F227",
	103 => X"D71F",
	104 => X"BE00",
	105 => X"A7F8",
	106 => X"960D",
	107 => X"8916",
	108 => X"81AE",
	109 => X"802F",
	110 => X"84A9",
	111 => X"8EE7",
	112 => X"9E70",
	113 => X"B288",
	114 => X"CA3F",
	115 => X"E47A",
	116 => X"0000",
	117 => X"1B83",
	118 => X"35BE",
	119 => X"4D75",
	120 => X"618D",
	121 => X"7116",
	122 => X"7B54",
	123 => X"7FCE",
	124 => X"7E4F",
	125 => X"76E7",
	126 => X"69F0",
	127 => X"5805",
	128 => X"41FD",
	129 => X"28DE",
	130 => X"0DD6",
	131 => X"F227",
	132 => X"D71F",
	133 => X"BE00",
	134 => X"A7F8",
	135 => X"960D",
	136 => X"8916",
	137 => X"81AE",
	138 => X"802F",
	139 => X"84A9",
	140 => X"8EE7",
	141 => X"9E70",
	142 => X"B288",
	143 => X"CA3F",
	144 => X"E47A",
	145 => X"0000",
	146 => X"1B83",
	147 => X"35BE",
	148 => X"4D75",
	149 => X"618D",
	150 => X"7116",
	151 => X"7B54",
	152 => X"7FCE",
	153 => X"7E4F",
	154 => X"76E7",
	155 => X"69F0",
	156 => X"5805",
	157 => X"41FD",
	158 => X"28DE",
	159 => X"0DD6",
	160 => X"F227",
	161 => X"D71F",
	162 => X"BE00",
	163 => X"A7F8",
	164 => X"960D",
	165 => X"8916",
	166 => X"81AE",
	167 => X"802F",
	168 => X"84A9",
	169 => X"8EE7",
	170 => X"9E70",
	171 => X"B288",
	172 => X"CA3F",
	173 => X"E47A",
	174 => X"0000",
	175 => X"1B83",
	176 => X"35BE",
	177 => X"4D75",
	178 => X"618D",
	179 => X"7116",
	180 => X"7B54",
	181 => X"7FCE",
	182 => X"7E4F",
	183 => X"76E7",
	184 => X"69F0",
	185 => X"5805",
	186 => X"41FD",
	187 => X"28DE",
	188 => X"0DD6",
	189 => X"F227",
	190 => X"D71F",
	191 => X"BE00",
	192 => X"A7F8",
	193 => X"960D",
	194 => X"8916",
	195 => X"81AE",
	196 => X"802F",
	197 => X"84A9",
	198 => X"8EE7",
	199 => X"9E70",
	200 => X"B288",
	201 => X"CA3F",
	202 => X"E47A",
	203 => X"0000",
	204 => X"1B83",
	205 => X"35BE",
	206 => X"4D75",
	207 => X"618D",
	208 => X"7116",
	209 => X"7B54",
	210 => X"7FCE",
	211 => X"7E4F",
	212 => X"76E7",
	213 => X"69F0",
	214 => X"5805",
	215 => X"41FD",
	216 => X"28DE",
	217 => X"0DD6",
	218 => X"F227",
	219 => X"D71F",
	220 => X"BE00",
	221 => X"A7F8",
	222 => X"960D",
	223 => X"8916",
	224 => X"81AE",
	225 => X"802F",
	226 => X"84A9",
	227 => X"8EE7",
	228 => X"9E70",
	229 => X"B288",
	230 => X"CA3F",
	231 => X"E47A",
	232 => X"0000",
	233 => X"1B83",
	234 => X"35BE",
	235 => X"4D75",
	236 => X"618D",
	237 => X"7116",
	238 => X"7B54",
	239 => X"7FCE",
	240 => X"7E4F",
	241 => X"76E7",
	242 => X"69F0",
	243 => X"5805",
	244 => X"41FD",
	245 => X"28DE",
	246 => X"0DD6",
	247 => X"F227",
	others => X"0000"
);

CONSTANT D6: hex := (
	000 => X"0000",
	001 => X"1C7B",
	002 => X"3789",
	003 => X"4FCD",
	004 => X"6412",
	005 => X"7352",
	006 => X"7CC9",
	007 => X"7FFF",
	008 => X"7CC9",
	009 => X"7352",
	010 => X"6412",
	011 => X"4FCD",
	012 => X"3789",
	013 => X"1C7B",
	014 => X"FFFD",
	015 => X"E382",
	016 => X"C874",
	017 => X"B030",
	018 => X"9BEB",
	019 => X"8CAB",
	020 => X"8334",
	021 => X"7FFF",
	022 => X"8334",
	023 => X"8CAB",
	024 => X"9BEB",
	025 => X"B030",
	026 => X"C874",
	027 => X"E382",
	028 => X"FFFD",
	029 => X"1C7B",
	030 => X"3789",
	031 => X"4FCD",
	032 => X"6412",
	033 => X"7352",
	034 => X"7CC9",
	035 => X"7FFF",
	036 => X"7CC9",
	037 => X"7352",
	038 => X"6412",
	039 => X"4FCD",
	040 => X"3789",
	041 => X"1C7B",
	042 => X"0000",
	043 => X"E382",
	044 => X"C874",
	045 => X"B030",
	046 => X"9BEB",
	047 => X"8CAB",
	048 => X"8334",
	049 => X"7FFF",
	050 => X"8334",
	051 => X"8CAB",
	052 => X"9BEB",
	053 => X"B030",
	054 => X"C874",
	055 => X"E382",
	056 => X"0000",
	057 => X"1C7B",
	058 => X"3789",
	059 => X"4FCD",
	060 => X"6412",
	061 => X"7352",
	062 => X"7CC9",
	063 => X"7FFF",
	064 => X"7CC9",
	065 => X"7352",
	066 => X"6412",
	067 => X"4FCD",
	068 => X"3789",
	069 => X"1C7B",
	070 => X"FFFD",
	071 => X"E382",
	072 => X"C874",
	073 => X"B030",
	074 => X"9BEB",
	075 => X"8CAB",
	076 => X"8334",
	077 => X"7FFF",
	078 => X"8334",
	079 => X"8CAB",
	080 => X"9BEB",
	081 => X"B030",
	082 => X"C874",
	083 => X"E382",
	084 => X"0000",
	085 => X"1C7B",
	086 => X"3789",
	087 => X"4FCD",
	088 => X"6412",
	089 => X"7352",
	090 => X"7CC9",
	091 => X"7FFF",
	092 => X"7CC9",
	093 => X"7352",
	094 => X"6412",
	095 => X"4FCD",
	096 => X"3789",
	097 => X"1C7B",
	098 => X"FFFD",
	099 => X"E382",
	100 => X"C874",
	101 => X"B030",
	102 => X"9BEB",
	103 => X"8CAB",
	104 => X"8334",
	105 => X"7FFF",
	106 => X"8334",
	107 => X"8CAB",
	108 => X"9BEB",
	109 => X"B030",
	110 => X"C874",
	111 => X"E382",
	112 => X"0000",
	113 => X"1C7B",
	114 => X"3789",
	115 => X"4FCD",
	116 => X"6412",
	117 => X"7352",
	118 => X"7CC9",
	119 => X"7FFF",
	120 => X"7CC9",
	121 => X"7352",
	122 => X"6412",
	123 => X"4FCD",
	124 => X"3789",
	125 => X"1C7B",
	126 => X"FFFD",
	127 => X"E382",
	128 => X"C874",
	129 => X"B030",
	130 => X"9BEB",
	131 => X"8CAB",
	132 => X"8334",
	133 => X"7FFF",
	134 => X"8334",
	135 => X"8CAB",
	136 => X"9BEB",
	137 => X"B030",
	138 => X"C874",
	139 => X"E382",
	140 => X"0000",
	141 => X"1C7B",
	142 => X"3789",
	143 => X"4FCD",
	144 => X"6412",
	145 => X"7352",
	146 => X"7CC9",
	147 => X"7FFF",
	148 => X"7CC9",
	149 => X"7352",
	150 => X"6412",
	151 => X"4FCD",
	152 => X"3789",
	153 => X"1C7B",
	154 => X"FFFD",
	155 => X"E382",
	156 => X"C874",
	157 => X"B030",
	158 => X"9BEB",
	159 => X"8CAB",
	160 => X"8334",
	161 => X"7FFF",
	162 => X"8334",
	163 => X"8CAB",
	164 => X"9BEB",
	165 => X"B030",
	166 => X"C874",
	167 => X"E382",
	168 => X"0000",
	169 => X"1C7B",
	170 => X"3789",
	171 => X"4FCD",
	172 => X"6412",
	173 => X"7352",
	174 => X"7CC9",
	175 => X"7FFF",
	176 => X"7CC9",
	177 => X"7352",
	178 => X"6412",
	179 => X"4FCD",
	180 => X"3789",
	181 => X"1C7B",
	182 => X"0000",
	183 => X"E382",
	184 => X"C874",
	185 => X"B030",
	186 => X"9BEB",
	187 => X"8CAB",
	188 => X"8334",
	189 => X"7FFF",
	190 => X"8334",
	191 => X"8CAB",
	192 => X"9BEB",
	193 => X"B030",
	194 => X"C874",
	195 => X"E382",
	196 => X"FFFD",
	197 => X"1C7B",
	198 => X"3789",
	199 => X"4FCD",
	200 => X"6412",
	201 => X"7352",
	202 => X"7CC9",
	203 => X"7FFF",
	204 => X"7CC9",
	205 => X"7352",
	206 => X"6412",
	207 => X"4FCD",
	208 => X"3789",
	209 => X"1C7B",
	210 => X"0000",
	211 => X"E382",
	212 => X"C874",
	213 => X"B030",
	214 => X"9BEB",
	215 => X"8CAB",
	216 => X"8334",
	217 => X"7FFF",
	218 => X"8334",
	219 => X"8CAB",
	220 => X"9BEB",
	221 => X"B030",
	222 => X"C874",
	223 => X"E382",
	224 => X"FFFD",
	225 => X"1C7B",
	226 => X"3789",
	227 => X"4FCD",
	228 => X"6412",
	229 => X"7352",
	230 => X"7CC9",
	231 => X"7FFF",
	232 => X"7CC9",
	233 => X"7352",
	234 => X"6412",
	235 => X"4FCD",
	236 => X"3789",
	237 => X"1C7B",
	238 => X"0000",
	239 => X"E382",
	240 => X"C874",
	241 => X"B030",
	242 => X"9BEB",
	243 => X"8CAB",
	244 => X"8334",
	245 => X"7FFF",
	246 => X"8334",
	247 => X"8CAB",
	others => X"0000"
);

CONSTANT DS6: hex := (
	000 => X"0000",
	001 => X"1EA1",
	002 => X"3B7B",
	003 => X"54E0",
	004 => X"6956",
	005 => X"77AD",
	006 => X"7F10",
	007 => X"7F10",
	008 => X"77AD",
	009 => X"6956",
	010 => X"54E0",
	011 => X"3B7B",
	012 => X"1EA1",
	013 => X"0000",
	014 => X"E15C",
	015 => X"C482",
	016 => X"AB1D",
	017 => X"96A7",
	018 => X"8850",
	019 => X"80ED",
	020 => X"80ED",
	021 => X"8850",
	022 => X"96A7",
	023 => X"AB1D",
	024 => X"C482",
	025 => X"E15C",
	026 => X"0000",
	027 => X"1EA1",
	028 => X"3B7B",
	029 => X"54E0",
	030 => X"6956",
	031 => X"77AD",
	032 => X"7F10",
	033 => X"7F10",
	034 => X"77AD",
	035 => X"6956",
	036 => X"54E0",
	037 => X"3B7B",
	038 => X"1EA1",
	039 => X"FFFD",
	040 => X"E15C",
	041 => X"C482",
	042 => X"AB1D",
	043 => X"96A7",
	044 => X"8850",
	045 => X"80ED",
	046 => X"80ED",
	047 => X"8850",
	048 => X"96A7",
	049 => X"AB1D",
	050 => X"C482",
	051 => X"E15C",
	052 => X"FFFD",
	053 => X"1EA1",
	054 => X"3B7B",
	055 => X"54E0",
	056 => X"6956",
	057 => X"77AD",
	058 => X"7F10",
	059 => X"7F10",
	060 => X"77AD",
	061 => X"6956",
	062 => X"54E0",
	063 => X"3B7B",
	064 => X"1EA1",
	065 => X"0000",
	066 => X"E15C",
	067 => X"C482",
	068 => X"AB1D",
	069 => X"96A7",
	070 => X"8850",
	071 => X"80ED",
	072 => X"80ED",
	073 => X"8850",
	074 => X"96A7",
	075 => X"AB1D",
	076 => X"C482",
	077 => X"E15C",
	078 => X"FFFD",
	079 => X"1EA1",
	080 => X"3B7B",
	081 => X"54E0",
	082 => X"6956",
	083 => X"77AD",
	084 => X"7F10",
	085 => X"7F10",
	086 => X"77AD",
	087 => X"6956",
	088 => X"54E0",
	089 => X"3B7B",
	090 => X"1EA1",
	091 => X"0000",
	092 => X"E15C",
	093 => X"C482",
	094 => X"AB1D",
	095 => X"96A7",
	096 => X"8850",
	097 => X"80ED",
	098 => X"80ED",
	099 => X"8850",
	100 => X"96A7",
	101 => X"AB1D",
	102 => X"C482",
	103 => X"E15C",
	104 => X"FFFD",
	105 => X"1EA1",
	106 => X"3B7B",
	107 => X"54E0",
	108 => X"6956",
	109 => X"77AD",
	110 => X"7F10",
	111 => X"7F10",
	112 => X"77AD",
	113 => X"6956",
	114 => X"54E0",
	115 => X"3B7B",
	116 => X"1EA1",
	117 => X"0000",
	118 => X"E15C",
	119 => X"C482",
	120 => X"AB1D",
	121 => X"96A7",
	122 => X"8850",
	123 => X"80ED",
	124 => X"80ED",
	125 => X"8850",
	126 => X"96A7",
	127 => X"AB1D",
	128 => X"C482",
	129 => X"E15C",
	130 => X"FFFD",
	131 => X"1EA1",
	132 => X"3B7B",
	133 => X"54E0",
	134 => X"6956",
	135 => X"77AD",
	136 => X"7F10",
	137 => X"7F10",
	138 => X"77AD",
	139 => X"6956",
	140 => X"54E0",
	141 => X"3B7B",
	142 => X"1EA1",
	143 => X"0000",
	144 => X"E15C",
	145 => X"C482",
	146 => X"AB1D",
	147 => X"96A7",
	148 => X"8850",
	149 => X"80ED",
	150 => X"80ED",
	151 => X"8850",
	152 => X"96A7",
	153 => X"AB1D",
	154 => X"C482",
	155 => X"E15C",
	156 => X"FFFD",
	157 => X"1EA1",
	158 => X"3B7B",
	159 => X"54E0",
	160 => X"6956",
	161 => X"77AD",
	162 => X"7F10",
	163 => X"7F10",
	164 => X"77AD",
	165 => X"6956",
	166 => X"54E0",
	167 => X"3B7B",
	168 => X"1EA1",
	169 => X"0000",
	170 => X"E15C",
	171 => X"C482",
	172 => X"AB1D",
	173 => X"96A7",
	174 => X"8850",
	175 => X"80ED",
	176 => X"80ED",
	177 => X"8850",
	178 => X"96A7",
	179 => X"AB1D",
	180 => X"C482",
	181 => X"E15C",
	182 => X"FFFD",
	183 => X"1EA1",
	184 => X"3B7B",
	185 => X"54E0",
	186 => X"6956",
	187 => X"77AD",
	188 => X"7F10",
	189 => X"7F10",
	190 => X"77AD",
	191 => X"6956",
	192 => X"54E0",
	193 => X"3B7B",
	194 => X"1EA1",
	195 => X"0000",
	196 => X"E15C",
	197 => X"C482",
	198 => X"AB1D",
	199 => X"96A7",
	200 => X"8850",
	201 => X"80ED",
	202 => X"80ED",
	203 => X"8850",
	204 => X"96A7",
	205 => X"AB1D",
	206 => X"C482",
	207 => X"E15C",
	208 => X"FFFD",
	209 => X"1EA1",
	210 => X"3B7B",
	211 => X"54E0",
	212 => X"6956",
	213 => X"77AD",
	214 => X"7F10",
	215 => X"7F10",
	216 => X"77AD",
	217 => X"6956",
	218 => X"54E0",
	219 => X"3B7B",
	220 => X"1EA1",
	221 => X"0000",
	222 => X"E15C",
	223 => X"C482",
	224 => X"AB1D",
	225 => X"96A7",
	226 => X"8850",
	227 => X"80ED",
	228 => X"80ED",
	229 => X"8850",
	230 => X"96A7",
	231 => X"AB1D",
	232 => X"C482",
	233 => X"E15C",
	234 => X"FFFD",
	235 => X"1EA1",
	236 => X"3B7B",
	237 => X"54E0",
	238 => X"6956",
	239 => X"77AD",
	240 => X"7F10",
	241 => X"7F10",
	242 => X"77AD",
	243 => X"6956",
	244 => X"54E0",
	245 => X"3B7B",
	246 => X"1EA1",
	247 => X"0000",
	others => X"0000"
);

BEGIN

--map all notes
key15_map: SampleContainer port map(clk, keys(15), C3, C4, C5, num_samples(015), num_samples(115), num_samples(215), octave, audio_request, k15);
key14_map: SampleContainer port map(clk, keys(14), CS3, CS4, CS5, num_samples(014), num_samples(114), num_samples(214), octave, audio_request, k14);
key13_map: SampleContainer port map(clk, keys(13), D3, D4, D5, num_samples(013), num_samples(113), num_samples(213), octave, audio_request, k13);
key12_map: SampleContainer port map(clk, keys(12), DS3, DS4, DS5, num_samples(012), num_samples(112), num_samples(212), octave, audio_request, k12);
key11_map: SampleContainer port map(clk, keys(11), E3, E4, E5, num_samples(011), num_samples(111), num_samples(211), octave, audio_request, k11);
key10_map: SampleContainer port map(clk, keys(10), F3, F4, F5, num_samples(010), num_samples(110), num_samples(210), octave, audio_request, k10);
--key9_map: SampleContainer port map(clk, keys(9), FS3, FS4, FS5, num_samples(009), num_samples(109), num_samples(209), octave, audio_request, k9);
--key8_map: SampleContainer port map(clk, keys(8), G3, G4, G5, num_samples(008), num_samples(108), num_samples(208), octave, audio_request, k8);
--key7_map: SampleContainer port map(clk, keys(7), GS3, GS4, GS5, num_samples(007), num_samples(107), num_samples(207), octave, audio_request, k7);
--key6_map: SampleContainer port map(clk, keys(6), A3, A4, A5, num_samples(006), num_samples(106), num_samples(206), octave, audio_request, k6);
--key5_map: SampleContainer port map(clk, keys(5), AS3, AS4, AS5, num_samples(005), num_samples(105), num_samples(205), octave, audio_request, k5);
--key4_map: SampleContainer port map(clk, keys(4), B3, B4, B5, num_samples(004), num_samples(104), num_samples(204), octave, audio_request, k4);
--key3_map: SampleContainer port map(clk, keys(3), C4, C5, C6, num_samples(003), num_samples(103), num_samples(203), octave, audio_request, k3);
--key2_map: SampleContainer port map(clk, keys(2), CS4, CS5, CS6, num_samples(002), num_samples(102), num_samples(202), octave, audio_request, k2);
--key1_map: SampleContainer port map(clk, keys(1), D4, D5, D6, num_samples(001), num_samples(101), num_samples(201), octave, audio_request, k1);
--key0_map: SampleContainer port map(clk, keys(0), DS4, DS5, DS6, num_samples(000), num_samples(100), num_samples(200), octave, audio_request, k0);

sample_adder: SampleAdder16 port map(keys, k0, k1, k2, k3, k4, k5, k6, k7, k8, k9, k10, k11, k12, k13, k14, k15, z);

END ARCHITECTURE rom;