library ieee;
use ieee.std_logic_1164.all;

package constants is
	constant DATA_SIZE : integer := 16;
	end package constants;
	
package body constants is
end package body constants;